module picorv32 (clk, resetn, mem_ready, mem_rdata, pcpi_wr, pcpi_rd, pcpi_wait, pcpi_ready, irq, trap, mem_valid, mem_instr, mem_addr, mem_wdata, mem_wstrb, mem_la_read, mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid, pcpi_insn, pcpi_rs1, pcpi_rs2, eoi, trace_valid, trace_data);

input clk;
input resetn;
input mem_ready;
input pcpi_wr;
input pcpi_wait;
input pcpi_ready;
output trap;
output mem_valid;
output mem_instr;
output mem_la_read;
output mem_la_write;
output pcpi_valid;
output trace_valid;
input [31:0] mem_rdata;
input [31:0] pcpi_rd;
input [31:0] irq;
output [31:0] mem_addr;
output [31:0] mem_wdata;
output [3:0] mem_wstrb;
output [31:0] mem_la_addr;
output [31:0] mem_la_wdata;
output [3:0] mem_la_wstrb;
output [31:0] pcpi_insn;
output [31:0] pcpi_rs1;
output [31:0] pcpi_rs2;
output [31:0] eoi;
output [35:0] trace_data;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(_7556_), .Y(_7556__hier0_bF_buf5) );
BUFX2 BUFX2_2 ( .A(_7556_), .Y(_7556__hier0_bF_buf4) );
BUFX2 BUFX2_3 ( .A(_7556_), .Y(_7556__hier0_bF_buf3) );
BUFX2 BUFX2_4 ( .A(_7556_), .Y(_7556__hier0_bF_buf2) );
BUFX2 BUFX2_5 ( .A(_7556_), .Y(_7556__hier0_bF_buf1) );
BUFX2 BUFX2_6 ( .A(_7556_), .Y(_7556__hier0_bF_buf0) );
BUFX2 BUFX2_7 ( .A(clk), .Y(clk_hier0_bF_buf10) );
BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf9) );
BUFX2 BUFX2_9 ( .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX2 BUFX2_10 ( .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX2 BUFX2_11 ( .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX2 BUFX2_12 ( .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX2 BUFX2_13 ( .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX2 BUFX2_14 ( .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX2 BUFX2_15 ( .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX2 BUFX2_16 ( .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX2 BUFX2_17 ( .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX2 BUFX2_18 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf5) );
BUFX2 BUFX2_19 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf4) );
BUFX2 BUFX2_20 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf3) );
BUFX2 BUFX2_21 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf2) );
BUFX2 BUFX2_22 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf1) );
BUFX2 BUFX2_23 ( .A(decoded_rs2_1_), .Y(decoded_rs2_1__hier0_bF_buf0) );
BUFX2 BUFX2_24 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf5) );
BUFX2 BUFX2_25 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf4) );
BUFX2 BUFX2_26 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf3) );
BUFX2 BUFX2_27 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf2) );
BUFX2 BUFX2_28 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf1) );
BUFX2 BUFX2_29 ( .A(decoded_rs1_1_), .Y(decoded_rs1_1__hier0_bF_buf0) );
BUFX2 BUFX2_30 ( .A(_7569_), .Y(_7569__hier0_bF_buf6) );
BUFX2 BUFX2_31 ( .A(_7569_), .Y(_7569__hier0_bF_buf5) );
BUFX2 BUFX2_32 ( .A(_7569_), .Y(_7569__hier0_bF_buf4) );
BUFX2 BUFX2_33 ( .A(_7569_), .Y(_7569__hier0_bF_buf3) );
BUFX2 BUFX2_34 ( .A(_7569_), .Y(_7569__hier0_bF_buf2) );
BUFX2 BUFX2_35 ( .A(_7569_), .Y(_7569__hier0_bF_buf1) );
BUFX2 BUFX2_36 ( .A(_7569_), .Y(_7569__hier0_bF_buf0) );
BUFX2 BUFX2_37 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf7) );
BUFX2 BUFX2_38 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf6) );
BUFX2 BUFX2_39 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf5) );
BUFX2 BUFX2_40 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf4) );
BUFX2 BUFX2_41 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf3) );
BUFX2 BUFX2_42 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf2) );
BUFX2 BUFX2_43 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf1) );
BUFX2 BUFX2_44 ( .A(decoded_rs2_0_), .Y(decoded_rs2_0__hier0_bF_buf0) );
BUFX2 BUFX2_45 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf6) );
BUFX2 BUFX2_46 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf5) );
BUFX2 BUFX2_47 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf4) );
BUFX2 BUFX2_48 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf3) );
BUFX2 BUFX2_49 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf2) );
BUFX2 BUFX2_50 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf1) );
BUFX2 BUFX2_51 ( .A(decoded_rs1_0_), .Y(decoded_rs1_0__hier0_bF_buf0) );
BUFX2 BUFX2_52 ( .A(_1601_), .Y(_1601__bF_buf4) );
BUFX2 BUFX2_53 ( .A(_1601_), .Y(_1601__bF_buf3) );
BUFX2 BUFX2_54 ( .A(_1601_), .Y(_1601__bF_buf2) );
BUFX2 BUFX2_55 ( .A(_1601_), .Y(_1601__bF_buf1) );
BUFX2 BUFX2_56 ( .A(_1601_), .Y(_1601__bF_buf0) );
BUFX2 BUFX2_57 ( .A(_10099_), .Y(_10099__bF_buf3) );
BUFX2 BUFX2_58 ( .A(_10099_), .Y(_10099__bF_buf2) );
BUFX2 BUFX2_59 ( .A(_10099_), .Y(_10099__bF_buf1) );
BUFX2 BUFX2_60 ( .A(_10099_), .Y(_10099__bF_buf0) );
BUFX2 BUFX2_61 ( .A(_4587_), .Y(_4587__bF_buf3) );
BUFX2 BUFX2_62 ( .A(_4587_), .Y(_4587__bF_buf2) );
BUFX2 BUFX2_63 ( .A(_4587_), .Y(_4587__bF_buf1) );
BUFX2 BUFX2_64 ( .A(_4587_), .Y(_4587__bF_buf0) );
BUFX2 BUFX2_65 ( .A(_5813_), .Y(_5813__bF_buf7) );
BUFX2 BUFX2_66 ( .A(_5813_), .Y(_5813__bF_buf6) );
BUFX2 BUFX2_67 ( .A(_5813_), .Y(_5813__bF_buf5) );
BUFX2 BUFX2_68 ( .A(_5813_), .Y(_5813__bF_buf4) );
BUFX2 BUFX2_69 ( .A(_5813_), .Y(_5813__bF_buf3) );
BUFX2 BUFX2_70 ( .A(_5813_), .Y(_5813__bF_buf2) );
BUFX2 BUFX2_71 ( .A(_5813_), .Y(_5813__bF_buf1) );
BUFX2 BUFX2_72 ( .A(_5813_), .Y(_5813__bF_buf0) );
BUFX2 BUFX2_73 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf42) );
BUFX2 BUFX2_74 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf41) );
BUFX2 BUFX2_75 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf40) );
BUFX2 BUFX2_76 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf39) );
BUFX2 BUFX2_77 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf38) );
BUFX2 BUFX2_78 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf37) );
BUFX2 BUFX2_79 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf36) );
BUFX2 BUFX2_80 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf35) );
BUFX2 BUFX2_81 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf34) );
BUFX2 BUFX2_82 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf33) );
BUFX2 BUFX2_83 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf32) );
BUFX2 BUFX2_84 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf31) );
BUFX2 BUFX2_85 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf30) );
BUFX2 BUFX2_86 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf29) );
BUFX2 BUFX2_87 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf28) );
BUFX2 BUFX2_88 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf27) );
BUFX2 BUFX2_89 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf26) );
BUFX2 BUFX2_90 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf25) );
BUFX2 BUFX2_91 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf24) );
BUFX2 BUFX2_92 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf23) );
BUFX2 BUFX2_93 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf22) );
BUFX2 BUFX2_94 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf21) );
BUFX2 BUFX2_95 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf20) );
BUFX2 BUFX2_96 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf19) );
BUFX2 BUFX2_97 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf18) );
BUFX2 BUFX2_98 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf17) );
BUFX2 BUFX2_99 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf16) );
BUFX2 BUFX2_100 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf15) );
BUFX2 BUFX2_101 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf14) );
BUFX2 BUFX2_102 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf13) );
BUFX2 BUFX2_103 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf12) );
BUFX2 BUFX2_104 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf11) );
BUFX2 BUFX2_105 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf10) );
BUFX2 BUFX2_106 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf9) );
BUFX2 BUFX2_107 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf8) );
BUFX2 BUFX2_108 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf7) );
BUFX2 BUFX2_109 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf6) );
BUFX2 BUFX2_110 ( .A(_7556__hier0_bF_buf4), .Y(_7556__bF_buf5) );
BUFX2 BUFX2_111 ( .A(_7556__hier0_bF_buf3), .Y(_7556__bF_buf4) );
BUFX2 BUFX2_112 ( .A(_7556__hier0_bF_buf2), .Y(_7556__bF_buf3) );
BUFX2 BUFX2_113 ( .A(_7556__hier0_bF_buf1), .Y(_7556__bF_buf2) );
BUFX2 BUFX2_114 ( .A(_7556__hier0_bF_buf0), .Y(_7556__bF_buf1) );
BUFX2 BUFX2_115 ( .A(_7556__hier0_bF_buf5), .Y(_7556__bF_buf0) );
BUFX2 BUFX2_116 ( .A(_4740_), .Y(_4740__bF_buf4) );
BUFX2 BUFX2_117 ( .A(_4740_), .Y(_4740__bF_buf3) );
BUFX2 BUFX2_118 ( .A(_4740_), .Y(_4740__bF_buf2) );
BUFX2 BUFX2_119 ( .A(_4740_), .Y(_4740__bF_buf1) );
BUFX2 BUFX2_120 ( .A(_4740_), .Y(_4740__bF_buf0) );
BUFX2 BUFX2_121 ( .A(_4605_), .Y(_4605__bF_buf5) );
BUFX2 BUFX2_122 ( .A(_4605_), .Y(_4605__bF_buf4) );
BUFX2 BUFX2_123 ( .A(_4605_), .Y(_4605__bF_buf3) );
BUFX2 BUFX2_124 ( .A(_4605_), .Y(_4605__bF_buf2) );
BUFX2 BUFX2_125 ( .A(_4605_), .Y(_4605__bF_buf1) );
BUFX2 BUFX2_126 ( .A(_4605_), .Y(_4605__bF_buf0) );
BUFX2 BUFX2_127 ( .A(_3914_), .Y(_3914__bF_buf4) );
BUFX2 BUFX2_128 ( .A(_3914_), .Y(_3914__bF_buf3) );
BUFX2 BUFX2_129 ( .A(_3914_), .Y(_3914__bF_buf2) );
BUFX2 BUFX2_130 ( .A(_3914_), .Y(_3914__bF_buf1) );
BUFX2 BUFX2_131 ( .A(_3914_), .Y(_3914__bF_buf0) );
BUFX2 BUFX2_132 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf8_) );
BUFX2 BUFX2_133 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf7_) );
BUFX2 BUFX2_134 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf6_) );
BUFX2 BUFX2_135 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf5_) );
BUFX2 BUFX2_136 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf4_) );
BUFX2 BUFX2_137 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf3_) );
BUFX2 BUFX2_138 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf2_) );
BUFX2 BUFX2_139 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf1_) );
BUFX2 BUFX2_140 ( .A(decoded_rs2_2_), .Y(decoded_rs2_2_bF_buf0_) );
BUFX2 BUFX2_141 ( .A(_2171_), .Y(_2171__bF_buf8) );
BUFX2 BUFX2_142 ( .A(_2171_), .Y(_2171__bF_buf7) );
BUFX2 BUFX2_143 ( .A(_2171_), .Y(_2171__bF_buf6) );
BUFX2 BUFX2_144 ( .A(_2171_), .Y(_2171__bF_buf5) );
BUFX2 BUFX2_145 ( .A(_2171_), .Y(_2171__bF_buf4) );
BUFX2 BUFX2_146 ( .A(_2171_), .Y(_2171__bF_buf3) );
BUFX2 BUFX2_147 ( .A(_2171_), .Y(_2171__bF_buf2) );
BUFX2 BUFX2_148 ( .A(_2171_), .Y(_2171__bF_buf1) );
BUFX2 BUFX2_149 ( .A(_2171_), .Y(_2171__bF_buf0) );
BUFX2 BUFX2_150 ( .A(_5140_), .Y(_5140__bF_buf5) );
BUFX2 BUFX2_151 ( .A(_5140_), .Y(_5140__bF_buf4) );
BUFX2 BUFX2_152 ( .A(_5140_), .Y(_5140__bF_buf3) );
BUFX2 BUFX2_153 ( .A(_5140_), .Y(_5140__bF_buf2) );
BUFX2 BUFX2_154 ( .A(_5140_), .Y(_5140__bF_buf1) );
BUFX2 BUFX2_155 ( .A(_5140_), .Y(_5140__bF_buf0) );
BUFX2 BUFX2_156 ( .A(_4925_), .Y(_4925__bF_buf4) );
BUFX2 BUFX2_157 ( .A(_4925_), .Y(_4925__bF_buf3) );
BUFX2 BUFX2_158 ( .A(_4925_), .Y(_4925__bF_buf2) );
BUFX2 BUFX2_159 ( .A(_4925_), .Y(_4925__bF_buf1) );
BUFX2 BUFX2_160 ( .A(_4925_), .Y(_4925__bF_buf0) );
BUFX2 BUFX2_161 ( .A(_4637_), .Y(_4637__bF_buf3) );
BUFX2 BUFX2_162 ( .A(_4637_), .Y(_4637__bF_buf2) );
BUFX2 BUFX2_163 ( .A(_4637_), .Y(_4637__bF_buf1) );
BUFX2 BUFX2_164 ( .A(_4637_), .Y(_4637__bF_buf0) );
BUFX2 BUFX2_165 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf12_) );
BUFX2 BUFX2_166 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf11_) );
BUFX2 BUFX2_167 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf10_) );
BUFX2 BUFX2_168 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf9_) );
BUFX2 BUFX2_169 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf8_) );
BUFX2 BUFX2_170 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf7_) );
BUFX2 BUFX2_171 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf6_) );
BUFX2 BUFX2_172 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf5_) );
BUFX2 BUFX2_173 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf4_) );
BUFX2 BUFX2_174 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf3_) );
BUFX2 BUFX2_175 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf2_) );
BUFX2 BUFX2_176 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf1_) );
BUFX2 BUFX2_177 ( .A(decoded_rs1_2_), .Y(decoded_rs1_2_bF_buf0_) );
BUFX2 BUFX2_178 ( .A(_3755_), .Y(_3755__bF_buf3) );
BUFX2 BUFX2_179 ( .A(_3755_), .Y(_3755__bF_buf2) );
BUFX2 BUFX2_180 ( .A(_3755_), .Y(_3755__bF_buf1) );
BUFX2 BUFX2_181 ( .A(_3755_), .Y(_3755__bF_buf0) );
BUFX2 BUFX2_182 ( .A(_1630_), .Y(_1630__bF_buf3) );
BUFX2 BUFX2_183 ( .A(_1630_), .Y(_1630__bF_buf2) );
BUFX2 BUFX2_184 ( .A(_1630_), .Y(_1630__bF_buf1) );
BUFX2 BUFX2_185 ( .A(_1630_), .Y(_1630__bF_buf0) );
BUFX2 BUFX2_186 ( .A(_2071_), .Y(_2071__bF_buf4) );
BUFX2 BUFX2_187 ( .A(_2071_), .Y(_2071__bF_buf3) );
BUFX2 BUFX2_188 ( .A(_2071_), .Y(_2071__bF_buf2) );
BUFX2 BUFX2_189 ( .A(_2071_), .Y(_2071__bF_buf1) );
BUFX2 BUFX2_190 ( .A(_2071_), .Y(_2071__bF_buf0) );
BUFX2 BUFX2_191 ( .A(cpu_state_5_), .Y(cpu_state_5_bF_buf3_) );
BUFX2 BUFX2_192 ( .A(cpu_state_5_), .Y(cpu_state_5_bF_buf2_) );
BUFX2 BUFX2_193 ( .A(cpu_state_5_), .Y(cpu_state_5_bF_buf1_) );
BUFX2 BUFX2_194 ( .A(cpu_state_5_), .Y(cpu_state_5_bF_buf0_) );
BUFX2 BUFX2_195 ( .A(_5707_), .Y(_5707__bF_buf3) );
BUFX2 BUFX2_196 ( .A(_5707_), .Y(_5707__bF_buf2) );
BUFX2 BUFX2_197 ( .A(_5707_), .Y(_5707__bF_buf1) );
BUFX2 BUFX2_198 ( .A(_5707_), .Y(_5707__bF_buf0) );
BUFX2 BUFX2_199 ( .A(_4731_), .Y(_4731__bF_buf4) );
BUFX2 BUFX2_200 ( .A(_4731_), .Y(_4731__bF_buf3) );
BUFX2 BUFX2_201 ( .A(_4731_), .Y(_4731__bF_buf2) );
BUFX2 BUFX2_202 ( .A(_4731_), .Y(_4731__bF_buf1) );
BUFX2 BUFX2_203 ( .A(_4731_), .Y(_4731__bF_buf0) );
BUFX2 BUFX2_204 ( .A(_4540_), .Y(_4540__bF_buf6) );
BUFX2 BUFX2_205 ( .A(_4540_), .Y(_4540__bF_buf5) );
BUFX2 BUFX2_206 ( .A(_4540_), .Y(_4540__bF_buf4) );
BUFX2 BUFX2_207 ( .A(_4540_), .Y(_4540__bF_buf3) );
BUFX2 BUFX2_208 ( .A(_4540_), .Y(_4540__bF_buf2) );
BUFX2 BUFX2_209 ( .A(_4540_), .Y(_4540__bF_buf1) );
BUFX2 BUFX2_210 ( .A(_4540_), .Y(_4540__bF_buf0) );
BUFX2 BUFX2_211 ( .A(_7700_), .Y(_7700__bF_buf5) );
BUFX2 BUFX2_212 ( .A(_7700_), .Y(_7700__bF_buf4) );
BUFX2 BUFX2_213 ( .A(_7700_), .Y(_7700__bF_buf3) );
BUFX2 BUFX2_214 ( .A(_7700_), .Y(_7700__bF_buf2) );
BUFX2 BUFX2_215 ( .A(_7700_), .Y(_7700__bF_buf1) );
BUFX2 BUFX2_216 ( .A(_7700_), .Y(_7700__bF_buf0) );
BUFX2 BUFX2_217 ( .A(_10728__3_), .Y(_10728__3_bF_buf4_) );
BUFX2 BUFX2_218 ( .A(_10728__3_), .Y(_10728__3_bF_buf3_) );
BUFX2 BUFX2_219 ( .A(_10728__3_), .Y(_10728__3_bF_buf2_) );
BUFX2 BUFX2_220 ( .A(_10728__3_), .Y(_10728__3_bF_buf1_) );
BUFX2 BUFX2_221 ( .A(_10728__3_), .Y(_10728__3_bF_buf0_) );
BUFX2 BUFX2_222 ( .A(_4863_), .Y(_4863__bF_buf4) );
BUFX2 BUFX2_223 ( .A(_4863_), .Y(_4863__bF_buf3) );
BUFX2 BUFX2_224 ( .A(_4863_), .Y(_4863__bF_buf2) );
BUFX2 BUFX2_225 ( .A(_4863_), .Y(_4863__bF_buf1) );
BUFX2 BUFX2_226 ( .A(_4863_), .Y(_4863__bF_buf0) );
BUFX2 BUFX2_227 ( .A(_4919_), .Y(_4919__bF_buf4) );
BUFX2 BUFX2_228 ( .A(_4919_), .Y(_4919__bF_buf3) );
BUFX2 BUFX2_229 ( .A(_4919_), .Y(_4919__bF_buf2) );
BUFX2 BUFX2_230 ( .A(_4919_), .Y(_4919__bF_buf1) );
BUFX2 BUFX2_231 ( .A(_4919_), .Y(_4919__bF_buf0) );
BUFX2 BUFX2_232 ( .A(_3981_), .Y(_3981__bF_buf4) );
BUFX2 BUFX2_233 ( .A(_3981_), .Y(_3981__bF_buf3) );
BUFX2 BUFX2_234 ( .A(_3981_), .Y(_3981__bF_buf2) );
BUFX2 BUFX2_235 ( .A(_3981_), .Y(_3981__bF_buf1) );
BUFX2 BUFX2_236 ( .A(_3981_), .Y(_3981__bF_buf0) );
BUFX2 BUFX2_237 ( .A(_4575_), .Y(_4575__bF_buf4) );
BUFX2 BUFX2_238 ( .A(_4575_), .Y(_4575__bF_buf3) );
BUFX2 BUFX2_239 ( .A(_4575_), .Y(_4575__bF_buf2) );
BUFX2 BUFX2_240 ( .A(_4575_), .Y(_4575__bF_buf1) );
BUFX2 BUFX2_241 ( .A(_4575_), .Y(_4575__bF_buf0) );
BUFX2 BUFX2_242 ( .A(_3846_), .Y(_3846__bF_buf4) );
BUFX2 BUFX2_243 ( .A(_3846_), .Y(_3846__bF_buf3) );
BUFX2 BUFX2_244 ( .A(_3846_), .Y(_3846__bF_buf2) );
BUFX2 BUFX2_245 ( .A(_3846_), .Y(_3846__bF_buf1) );
BUFX2 BUFX2_246 ( .A(_3846_), .Y(_3846__bF_buf0) );
BUFX2 BUFX2_247 ( .A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4) );
BUFX2 BUFX2_248 ( .A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3) );
BUFX2 BUFX2_249 ( .A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2) );
BUFX2 BUFX2_250 ( .A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1) );
BUFX2 BUFX2_251 ( .A(is_lui_auipc_jal_jalr_addi_add_sub), .Y(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0) );
BUFX2 BUFX2_252 ( .A(latched_stalu), .Y(latched_stalu_bF_buf6) );
BUFX2 BUFX2_253 ( .A(latched_stalu), .Y(latched_stalu_bF_buf5) );
BUFX2 BUFX2_254 ( .A(latched_stalu), .Y(latched_stalu_bF_buf4) );
BUFX2 BUFX2_255 ( .A(latched_stalu), .Y(latched_stalu_bF_buf3) );
BUFX2 BUFX2_256 ( .A(latched_stalu), .Y(latched_stalu_bF_buf2) );
BUFX2 BUFX2_257 ( .A(latched_stalu), .Y(latched_stalu_bF_buf1) );
BUFX2 BUFX2_258 ( .A(latched_stalu), .Y(latched_stalu_bF_buf0) );
BUFX2 BUFX2_259 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf5_) );
BUFX2 BUFX2_260 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf4_) );
BUFX2 BUFX2_261 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf3_) );
BUFX2 BUFX2_262 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf2_) );
BUFX2 BUFX2_263 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf1_) );
BUFX2 BUFX2_264 ( .A(cpu_state_2_), .Y(cpu_state_2_bF_buf0_) );
BUFX2 BUFX2_265 ( .A(_1853_), .Y(_1853__bF_buf5) );
BUFX2 BUFX2_266 ( .A(_1853_), .Y(_1853__bF_buf4) );
BUFX2 BUFX2_267 ( .A(_1853_), .Y(_1853__bF_buf3) );
BUFX2 BUFX2_268 ( .A(_1853_), .Y(_1853__bF_buf2) );
BUFX2 BUFX2_269 ( .A(_1853_), .Y(_1853__bF_buf1) );
BUFX2 BUFX2_270 ( .A(_1853_), .Y(_1853__bF_buf0) );
BUFX2 BUFX2_271 ( .A(_5131_), .Y(_5131__bF_buf5) );
BUFX2 BUFX2_272 ( .A(_5131_), .Y(_5131__bF_buf4) );
BUFX2 BUFX2_273 ( .A(_5131_), .Y(_5131__bF_buf3) );
BUFX2 BUFX2_274 ( .A(_5131_), .Y(_5131__bF_buf2) );
BUFX2 BUFX2_275 ( .A(_5131_), .Y(_5131__bF_buf1) );
BUFX2 BUFX2_276 ( .A(_5131_), .Y(_5131__bF_buf0) );
BUFX2 BUFX2_277 ( .A(_5780_), .Y(_5780__bF_buf7) );
BUFX2 BUFX2_278 ( .A(_5780_), .Y(_5780__bF_buf6) );
BUFX2 BUFX2_279 ( .A(_5780_), .Y(_5780__bF_buf5) );
BUFX2 BUFX2_280 ( .A(_5780_), .Y(_5780__bF_buf4) );
BUFX2 BUFX2_281 ( .A(_5780_), .Y(_5780__bF_buf3) );
BUFX2 BUFX2_282 ( .A(_5780_), .Y(_5780__bF_buf2) );
BUFX2 BUFX2_283 ( .A(_5780_), .Y(_5780__bF_buf1) );
BUFX2 BUFX2_284 ( .A(_5780_), .Y(_5780__bF_buf0) );
BUFX2 BUFX2_285 ( .A(_10728__0_), .Y(_10728__0_bF_buf7_) );
BUFX2 BUFX2_286 ( .A(_10728__0_), .Y(_10728__0_bF_buf6_) );
BUFX2 BUFX2_287 ( .A(_10728__0_), .Y(_10728__0_bF_buf5_) );
BUFX2 BUFX2_288 ( .A(_10728__0_), .Y(_10728__0_bF_buf4_) );
BUFX2 BUFX2_289 ( .A(_10728__0_), .Y(_10728__0_bF_buf3_) );
BUFX2 BUFX2_290 ( .A(_10728__0_), .Y(_10728__0_bF_buf2_) );
BUFX2 BUFX2_291 ( .A(_10728__0_), .Y(_10728__0_bF_buf1_) );
BUFX2 BUFX2_292 ( .A(_10728__0_), .Y(_10728__0_bF_buf0_) );
BUFX2 BUFX2_293 ( .A(_3711_), .Y(_3711__bF_buf7) );
BUFX2 BUFX2_294 ( .A(_3711_), .Y(_3711__bF_buf6) );
BUFX2 BUFX2_295 ( .A(_3711_), .Y(_3711__bF_buf5) );
BUFX2 BUFX2_296 ( .A(_3711_), .Y(_3711__bF_buf4) );
BUFX2 BUFX2_297 ( .A(_3711_), .Y(_3711__bF_buf3) );
BUFX2 BUFX2_298 ( .A(_3711_), .Y(_3711__bF_buf2) );
BUFX2 BUFX2_299 ( .A(_3711_), .Y(_3711__bF_buf1) );
BUFX2 BUFX2_300 ( .A(_3711_), .Y(_3711__bF_buf0) );
BUFX2 BUFX2_301 ( .A(_4763_), .Y(_4763__bF_buf4) );
BUFX2 BUFX2_302 ( .A(_4763_), .Y(_4763__bF_buf3) );
BUFX2 BUFX2_303 ( .A(_4763_), .Y(_4763__bF_buf2) );
BUFX2 BUFX2_304 ( .A(_4763_), .Y(_4763__bF_buf1) );
BUFX2 BUFX2_305 ( .A(_4763_), .Y(_4763__bF_buf0) );
BUFX2 BUFX2_306 ( .A(decoder_trigger), .Y(decoder_trigger_bF_buf3) );
BUFX2 BUFX2_307 ( .A(decoder_trigger), .Y(decoder_trigger_bF_buf2) );
BUFX2 BUFX2_308 ( .A(decoder_trigger), .Y(decoder_trigger_bF_buf1) );
BUFX2 BUFX2_309 ( .A(decoder_trigger), .Y(decoder_trigger_bF_buf0) );
BUFX2 BUFX2_310 ( .A(instr_rdinstr), .Y(instr_rdinstr_bF_buf4) );
BUFX2 BUFX2_311 ( .A(instr_rdinstr), .Y(instr_rdinstr_bF_buf3) );
BUFX2 BUFX2_312 ( .A(instr_rdinstr), .Y(instr_rdinstr_bF_buf2) );
BUFX2 BUFX2_313 ( .A(instr_rdinstr), .Y(instr_rdinstr_bF_buf1) );
BUFX2 BUFX2_314 ( .A(instr_rdinstr), .Y(instr_rdinstr_bF_buf0) );
BUFX2 BUFX2_315 ( .A(_3746_), .Y(_3746__bF_buf3) );
BUFX2 BUFX2_316 ( .A(_3746_), .Y(_3746__bF_buf2) );
BUFX2 BUFX2_317 ( .A(_3746_), .Y(_3746__bF_buf1) );
BUFX2 BUFX2_318 ( .A(_3746_), .Y(_3746__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf136) );
CLKBUF1 CLKBUF1_2 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf135) );
CLKBUF1 CLKBUF1_3 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf134) );
CLKBUF1 CLKBUF1_4 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf133) );
CLKBUF1 CLKBUF1_5 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf132) );
CLKBUF1 CLKBUF1_6 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf131) );
CLKBUF1 CLKBUF1_7 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf130) );
CLKBUF1 CLKBUF1_8 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf129) );
CLKBUF1 CLKBUF1_9 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf128) );
CLKBUF1 CLKBUF1_10 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf127) );
CLKBUF1 CLKBUF1_11 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf126) );
CLKBUF1 CLKBUF1_12 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf125) );
CLKBUF1 CLKBUF1_13 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf124) );
CLKBUF1 CLKBUF1_14 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf123) );
CLKBUF1 CLKBUF1_15 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf122) );
CLKBUF1 CLKBUF1_16 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf121) );
CLKBUF1 CLKBUF1_17 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf120) );
CLKBUF1 CLKBUF1_18 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf119) );
CLKBUF1 CLKBUF1_19 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf118) );
CLKBUF1 CLKBUF1_20 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf117) );
CLKBUF1 CLKBUF1_21 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf116) );
CLKBUF1 CLKBUF1_22 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf115) );
CLKBUF1 CLKBUF1_23 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf114) );
CLKBUF1 CLKBUF1_24 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf113) );
CLKBUF1 CLKBUF1_25 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf112) );
CLKBUF1 CLKBUF1_26 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf111) );
CLKBUF1 CLKBUF1_27 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf110) );
CLKBUF1 CLKBUF1_28 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf109) );
CLKBUF1 CLKBUF1_29 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf108) );
CLKBUF1 CLKBUF1_30 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf107) );
CLKBUF1 CLKBUF1_31 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf106) );
CLKBUF1 CLKBUF1_32 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf105) );
CLKBUF1 CLKBUF1_33 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf104) );
CLKBUF1 CLKBUF1_34 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf103) );
CLKBUF1 CLKBUF1_35 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf102) );
CLKBUF1 CLKBUF1_36 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf101) );
CLKBUF1 CLKBUF1_37 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf100) );
CLKBUF1 CLKBUF1_38 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf99) );
CLKBUF1 CLKBUF1_39 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf98) );
CLKBUF1 CLKBUF1_40 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf97) );
CLKBUF1 CLKBUF1_41 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf96) );
CLKBUF1 CLKBUF1_42 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf95) );
CLKBUF1 CLKBUF1_43 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf94) );
CLKBUF1 CLKBUF1_44 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf93) );
CLKBUF1 CLKBUF1_45 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf92) );
CLKBUF1 CLKBUF1_46 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf91) );
CLKBUF1 CLKBUF1_47 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf90) );
CLKBUF1 CLKBUF1_48 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf89) );
CLKBUF1 CLKBUF1_49 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf88) );
CLKBUF1 CLKBUF1_50 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf87) );
CLKBUF1 CLKBUF1_51 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf86) );
CLKBUF1 CLKBUF1_52 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf85) );
CLKBUF1 CLKBUF1_53 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf84) );
CLKBUF1 CLKBUF1_54 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf83) );
CLKBUF1 CLKBUF1_55 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf82) );
CLKBUF1 CLKBUF1_56 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf81) );
CLKBUF1 CLKBUF1_57 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf80) );
CLKBUF1 CLKBUF1_58 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf79) );
CLKBUF1 CLKBUF1_59 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf78) );
CLKBUF1 CLKBUF1_60 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf77) );
CLKBUF1 CLKBUF1_61 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf76) );
CLKBUF1 CLKBUF1_62 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf75) );
CLKBUF1 CLKBUF1_63 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf74) );
CLKBUF1 CLKBUF1_64 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf73) );
CLKBUF1 CLKBUF1_65 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf72) );
CLKBUF1 CLKBUF1_66 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf71) );
CLKBUF1 CLKBUF1_67 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf70) );
CLKBUF1 CLKBUF1_68 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf69) );
CLKBUF1 CLKBUF1_69 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf68) );
CLKBUF1 CLKBUF1_70 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf67) );
CLKBUF1 CLKBUF1_71 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf66) );
CLKBUF1 CLKBUF1_72 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf65) );
CLKBUF1 CLKBUF1_73 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf64) );
CLKBUF1 CLKBUF1_74 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf63) );
CLKBUF1 CLKBUF1_75 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf62) );
CLKBUF1 CLKBUF1_76 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf61) );
CLKBUF1 CLKBUF1_77 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf60) );
CLKBUF1 CLKBUF1_78 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf59) );
CLKBUF1 CLKBUF1_79 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf58) );
CLKBUF1 CLKBUF1_80 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf57) );
CLKBUF1 CLKBUF1_81 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf56) );
CLKBUF1 CLKBUF1_82 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf55) );
CLKBUF1 CLKBUF1_83 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf54) );
CLKBUF1 CLKBUF1_84 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf53) );
CLKBUF1 CLKBUF1_85 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf52) );
CLKBUF1 CLKBUF1_86 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf51) );
CLKBUF1 CLKBUF1_87 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf50) );
CLKBUF1 CLKBUF1_88 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf49) );
CLKBUF1 CLKBUF1_89 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf48) );
CLKBUF1 CLKBUF1_90 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf47) );
CLKBUF1 CLKBUF1_91 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf46) );
CLKBUF1 CLKBUF1_92 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf45) );
CLKBUF1 CLKBUF1_93 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf44) );
CLKBUF1 CLKBUF1_94 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf43) );
CLKBUF1 CLKBUF1_95 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf42) );
CLKBUF1 CLKBUF1_96 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf41) );
CLKBUF1 CLKBUF1_97 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf40) );
CLKBUF1 CLKBUF1_98 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf39) );
CLKBUF1 CLKBUF1_99 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf38) );
CLKBUF1 CLKBUF1_100 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf37) );
CLKBUF1 CLKBUF1_101 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf36) );
CLKBUF1 CLKBUF1_102 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35) );
CLKBUF1 CLKBUF1_103 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf34) );
CLKBUF1 CLKBUF1_104 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf33) );
CLKBUF1 CLKBUF1_105 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf32) );
CLKBUF1 CLKBUF1_106 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf31) );
CLKBUF1 CLKBUF1_107 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf30) );
CLKBUF1 CLKBUF1_108 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf29) );
CLKBUF1 CLKBUF1_109 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
CLKBUF1 CLKBUF1_110 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf27) );
CLKBUF1 CLKBUF1_111 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf26) );
CLKBUF1 CLKBUF1_112 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf25) );
CLKBUF1 CLKBUF1_113 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf24) );
CLKBUF1 CLKBUF1_114 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf23) );
CLKBUF1 CLKBUF1_115 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf22) );
CLKBUF1 CLKBUF1_116 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf21) );
CLKBUF1 CLKBUF1_117 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf20) );
CLKBUF1 CLKBUF1_118 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf19) );
CLKBUF1 CLKBUF1_119 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf18) );
CLKBUF1 CLKBUF1_120 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf17) );
CLKBUF1 CLKBUF1_121 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf16) );
CLKBUF1 CLKBUF1_122 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf15) );
CLKBUF1 CLKBUF1_123 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf14) );
CLKBUF1 CLKBUF1_124 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf13) );
CLKBUF1 CLKBUF1_125 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf12) );
CLKBUF1 CLKBUF1_126 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_127 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_128 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_129 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_130 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_131 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_132 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_133 ( .A(clk_hier0_bF_buf10), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_134 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_135 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_136 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_137 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf0) );
BUFX2 BUFX2_319 ( .A(_4913_), .Y(_4913__bF_buf6) );
BUFX2 BUFX2_320 ( .A(_4913_), .Y(_4913__bF_buf5) );
BUFX2 BUFX2_321 ( .A(_4913_), .Y(_4913__bF_buf4) );
BUFX2 BUFX2_322 ( .A(_4913_), .Y(_4913__bF_buf3) );
BUFX2 BUFX2_323 ( .A(_4913_), .Y(_4913__bF_buf2) );
BUFX2 BUFX2_324 ( .A(_4913_), .Y(_4913__bF_buf1) );
BUFX2 BUFX2_325 ( .A(_4913_), .Y(_4913__bF_buf0) );
BUFX2 BUFX2_326 ( .A(_4722_), .Y(_4722__bF_buf4) );
BUFX2 BUFX2_327 ( .A(_4722_), .Y(_4722__bF_buf3) );
BUFX2 BUFX2_328 ( .A(_4722_), .Y(_4722__bF_buf2) );
BUFX2 BUFX2_329 ( .A(_4722_), .Y(_4722__bF_buf1) );
BUFX2 BUFX2_330 ( .A(_4722_), .Y(_4722__bF_buf0) );
BUFX2 BUFX2_331 ( .A(_4531_), .Y(_4531__bF_buf4) );
BUFX2 BUFX2_332 ( .A(_4531_), .Y(_4531__bF_buf3) );
BUFX2 BUFX2_333 ( .A(_4531_), .Y(_4531__bF_buf2) );
BUFX2 BUFX2_334 ( .A(_4531_), .Y(_4531__bF_buf1) );
BUFX2 BUFX2_335 ( .A(_4531_), .Y(_4531__bF_buf0) );
BUFX2 BUFX2_336 ( .A(_4816_), .Y(_4816__bF_buf4) );
BUFX2 BUFX2_337 ( .A(_4816_), .Y(_4816__bF_buf3) );
BUFX2 BUFX2_338 ( .A(_4816_), .Y(_4816__bF_buf2) );
BUFX2 BUFX2_339 ( .A(_4816_), .Y(_4816__bF_buf1) );
BUFX2 BUFX2_340 ( .A(_4816_), .Y(_4816__bF_buf0) );
BUFX2 BUFX2_341 ( .A(_4854_), .Y(_4854__bF_buf4) );
BUFX2 BUFX2_342 ( .A(_4854_), .Y(_4854__bF_buf3) );
BUFX2 BUFX2_343 ( .A(_4854_), .Y(_4854__bF_buf2) );
BUFX2 BUFX2_344 ( .A(_4854_), .Y(_4854__bF_buf1) );
BUFX2 BUFX2_345 ( .A(_4854_), .Y(_4854__bF_buf0) );
BUFX2 BUFX2_346 ( .A(_4014_), .Y(_4014__bF_buf7) );
BUFX2 BUFX2_347 ( .A(_4014_), .Y(_4014__bF_buf6) );
BUFX2 BUFX2_348 ( .A(_4014_), .Y(_4014__bF_buf5) );
BUFX2 BUFX2_349 ( .A(_4014_), .Y(_4014__bF_buf4) );
BUFX2 BUFX2_350 ( .A(_4014_), .Y(_4014__bF_buf3) );
BUFX2 BUFX2_351 ( .A(_4014_), .Y(_4014__bF_buf2) );
BUFX2 BUFX2_352 ( .A(_4014_), .Y(_4014__bF_buf1) );
BUFX2 BUFX2_353 ( .A(_4014_), .Y(_4014__bF_buf0) );
BUFX2 BUFX2_354 ( .A(_4948_), .Y(_4948__bF_buf4) );
BUFX2 BUFX2_355 ( .A(_4948_), .Y(_4948__bF_buf3) );
BUFX2 BUFX2_356 ( .A(_4948_), .Y(_4948__bF_buf2) );
BUFX2 BUFX2_357 ( .A(_4948_), .Y(_4948__bF_buf1) );
BUFX2 BUFX2_358 ( .A(_4948_), .Y(_4948__bF_buf0) );
BUFX2 BUFX2_359 ( .A(_7632_), .Y(_7632__bF_buf3) );
BUFX2 BUFX2_360 ( .A(_7632_), .Y(_7632__bF_buf2) );
BUFX2 BUFX2_361 ( .A(_7632_), .Y(_7632__bF_buf1) );
BUFX2 BUFX2_362 ( .A(_7632_), .Y(_7632__bF_buf0) );
BUFX2 BUFX2_363 ( .A(_7629_), .Y(_7629__bF_buf3) );
BUFX2 BUFX2_364 ( .A(_7629_), .Y(_7629__bF_buf2) );
BUFX2 BUFX2_365 ( .A(_7629_), .Y(_7629__bF_buf1) );
BUFX2 BUFX2_366 ( .A(_7629_), .Y(_7629__bF_buf0) );
BUFX2 BUFX2_367 ( .A(_4910_), .Y(_4910__bF_buf4) );
BUFX2 BUFX2_368 ( .A(_4910_), .Y(_4910__bF_buf3) );
BUFX2 BUFX2_369 ( .A(_4910_), .Y(_4910__bF_buf2) );
BUFX2 BUFX2_370 ( .A(_4910_), .Y(_4910__bF_buf1) );
BUFX2 BUFX2_371 ( .A(_4910_), .Y(_4910__bF_buf0) );
BUFX2 BUFX2_372 ( .A(_4431_), .Y(_4431__bF_buf7) );
BUFX2 BUFX2_373 ( .A(_4431_), .Y(_4431__bF_buf6) );
BUFX2 BUFX2_374 ( .A(_4431_), .Y(_4431__bF_buf5) );
BUFX2 BUFX2_375 ( .A(_4431_), .Y(_4431__bF_buf4) );
BUFX2 BUFX2_376 ( .A(_4431_), .Y(_4431__bF_buf3) );
BUFX2 BUFX2_377 ( .A(_4431_), .Y(_4431__bF_buf2) );
BUFX2 BUFX2_378 ( .A(_4431_), .Y(_4431__bF_buf1) );
BUFX2 BUFX2_379 ( .A(_4431_), .Y(_4431__bF_buf0) );
BUFX2 BUFX2_380 ( .A(_5348_), .Y(_5348__bF_buf5) );
BUFX2 BUFX2_381 ( .A(_5348_), .Y(_5348__bF_buf4) );
BUFX2 BUFX2_382 ( .A(_5348_), .Y(_5348__bF_buf3) );
BUFX2 BUFX2_383 ( .A(_5348_), .Y(_5348__bF_buf2) );
BUFX2 BUFX2_384 ( .A(_5348_), .Y(_5348__bF_buf1) );
BUFX2 BUFX2_385 ( .A(_5348_), .Y(_5348__bF_buf0) );
BUFX2 BUFX2_386 ( .A(_3223_), .Y(_3223__bF_buf3) );
BUFX2 BUFX2_387 ( .A(_3223_), .Y(_3223__bF_buf2) );
BUFX2 BUFX2_388 ( .A(_3223_), .Y(_3223__bF_buf1) );
BUFX2 BUFX2_389 ( .A(_3223_), .Y(_3223__bF_buf0) );
BUFX2 BUFX2_390 ( .A(_4713_), .Y(_4713__bF_buf4) );
BUFX2 BUFX2_391 ( .A(_4713_), .Y(_4713__bF_buf3) );
BUFX2 BUFX2_392 ( .A(_4713_), .Y(_4713__bF_buf2) );
BUFX2 BUFX2_393 ( .A(_4713_), .Y(_4713__bF_buf1) );
BUFX2 BUFX2_394 ( .A(_4713_), .Y(_4713__bF_buf0) );
BUFX2 BUFX2_395 ( .A(_4845_), .Y(_4845__bF_buf4) );
BUFX2 BUFX2_396 ( .A(_4845_), .Y(_4845__bF_buf3) );
BUFX2 BUFX2_397 ( .A(_4845_), .Y(_4845__bF_buf2) );
BUFX2 BUFX2_398 ( .A(_4845_), .Y(_4845__bF_buf1) );
BUFX2 BUFX2_399 ( .A(_4845_), .Y(_4845__bF_buf0) );
BUFX2 BUFX2_400 ( .A(_4654_), .Y(_4654__bF_buf4) );
BUFX2 BUFX2_401 ( .A(_4654_), .Y(_4654__bF_buf3) );
BUFX2 BUFX2_402 ( .A(_4654_), .Y(_4654__bF_buf2) );
BUFX2 BUFX2_403 ( .A(_4654_), .Y(_4654__bF_buf1) );
BUFX2 BUFX2_404 ( .A(_4654_), .Y(_4654__bF_buf0) );
BUFX2 BUFX2_405 ( .A(_5859_), .Y(_5859__bF_buf4) );
BUFX2 BUFX2_406 ( .A(_5859_), .Y(_5859__bF_buf3) );
BUFX2 BUFX2_407 ( .A(_5859_), .Y(_5859__bF_buf2) );
BUFX2 BUFX2_408 ( .A(_5859_), .Y(_5859__bF_buf1) );
BUFX2 BUFX2_409 ( .A(_5859_), .Y(_5859__bF_buf0) );
BUFX2 BUFX2_410 ( .A(_7623_), .Y(_7623__bF_buf4) );
BUFX2 BUFX2_411 ( .A(_7623_), .Y(_7623__bF_buf3) );
BUFX2 BUFX2_412 ( .A(_7623_), .Y(_7623__bF_buf2) );
BUFX2 BUFX2_413 ( .A(_7623_), .Y(_7623__bF_buf1) );
BUFX2 BUFX2_414 ( .A(_7623_), .Y(_7623__bF_buf0) );
BUFX2 BUFX2_415 ( .A(_4901_), .Y(_4901__bF_buf4) );
BUFX2 BUFX2_416 ( .A(_4901_), .Y(_4901__bF_buf3) );
BUFX2 BUFX2_417 ( .A(_4901_), .Y(_4901__bF_buf2) );
BUFX2 BUFX2_418 ( .A(_4901_), .Y(_4901__bF_buf1) );
BUFX2 BUFX2_419 ( .A(_4901_), .Y(_4901__bF_buf0) );
BUFX2 BUFX2_420 ( .A(_1967_), .Y(_1967__bF_buf6) );
BUFX2 BUFX2_421 ( .A(_1967_), .Y(_1967__bF_buf5) );
BUFX2 BUFX2_422 ( .A(_1967_), .Y(_1967__bF_buf4) );
BUFX2 BUFX2_423 ( .A(_1967_), .Y(_1967__bF_buf3) );
BUFX2 BUFX2_424 ( .A(_1967_), .Y(_1967__bF_buf2) );
BUFX2 BUFX2_425 ( .A(_1967_), .Y(_1967__bF_buf1) );
BUFX2 BUFX2_426 ( .A(_1967_), .Y(_1967__bF_buf0) );
BUFX2 BUFX2_427 ( .A(_1547_), .Y(_1547__bF_buf5) );
BUFX2 BUFX2_428 ( .A(_1547_), .Y(_1547__bF_buf4) );
BUFX2 BUFX2_429 ( .A(_1547_), .Y(_1547__bF_buf3) );
BUFX2 BUFX2_430 ( .A(_1547_), .Y(_1547__bF_buf2) );
BUFX2 BUFX2_431 ( .A(_1547_), .Y(_1547__bF_buf1) );
BUFX2 BUFX2_432 ( .A(_1547_), .Y(_1547__bF_buf0) );
BUFX2 BUFX2_433 ( .A(_5856_), .Y(_5856__bF_buf4) );
BUFX2 BUFX2_434 ( .A(_5856_), .Y(_5856__bF_buf3) );
BUFX2 BUFX2_435 ( .A(_5856_), .Y(_5856__bF_buf2) );
BUFX2 BUFX2_436 ( .A(_5856_), .Y(_5856__bF_buf1) );
BUFX2 BUFX2_437 ( .A(_5856_), .Y(_5856__bF_buf0) );
BUFX2 BUFX2_438 ( .A(_4783_), .Y(_4783__bF_buf4) );
BUFX2 BUFX2_439 ( .A(_4783_), .Y(_4783__bF_buf3) );
BUFX2 BUFX2_440 ( .A(_4783_), .Y(_4783__bF_buf2) );
BUFX2 BUFX2_441 ( .A(_4783_), .Y(_4783__bF_buf1) );
BUFX2 BUFX2_442 ( .A(_4783_), .Y(_4783__bF_buf0) );
BUFX2 BUFX2_443 ( .A(_7561_), .Y(_7561__bF_buf6) );
BUFX2 BUFX2_444 ( .A(_7561_), .Y(_7561__bF_buf5) );
BUFX2 BUFX2_445 ( .A(_7561_), .Y(_7561__bF_buf4) );
BUFX2 BUFX2_446 ( .A(_7561_), .Y(_7561__bF_buf3) );
BUFX2 BUFX2_447 ( .A(_7561_), .Y(_7561__bF_buf2) );
BUFX2 BUFX2_448 ( .A(_7561_), .Y(_7561__bF_buf1) );
BUFX2 BUFX2_449 ( .A(_7561_), .Y(_7561__bF_buf0) );
BUFX2 BUFX2_450 ( .A(_2138_), .Y(_2138__bF_buf4) );
BUFX2 BUFX2_451 ( .A(_2138_), .Y(_2138__bF_buf3) );
BUFX2 BUFX2_452 ( .A(_2138_), .Y(_2138__bF_buf2) );
BUFX2 BUFX2_453 ( .A(_2138_), .Y(_2138__bF_buf1) );
BUFX2 BUFX2_454 ( .A(_2138_), .Y(_2138__bF_buf0) );
BUFX2 BUFX2_455 ( .A(_4933_), .Y(_4933__bF_buf4) );
BUFX2 BUFX2_456 ( .A(_4933_), .Y(_4933__bF_buf3) );
BUFX2 BUFX2_457 ( .A(_4933_), .Y(_4933__bF_buf2) );
BUFX2 BUFX2_458 ( .A(_4933_), .Y(_4933__bF_buf1) );
BUFX2 BUFX2_459 ( .A(_4933_), .Y(_4933__bF_buf0) );
BUFX2 BUFX2_460 ( .A(instr_jal), .Y(instr_jal_bF_buf6) );
BUFX2 BUFX2_461 ( .A(instr_jal), .Y(instr_jal_bF_buf5) );
BUFX2 BUFX2_462 ( .A(instr_jal), .Y(instr_jal_bF_buf4) );
BUFX2 BUFX2_463 ( .A(instr_jal), .Y(instr_jal_bF_buf3) );
BUFX2 BUFX2_464 ( .A(instr_jal), .Y(instr_jal_bF_buf2) );
BUFX2 BUFX2_465 ( .A(instr_jal), .Y(instr_jal_bF_buf1) );
BUFX2 BUFX2_466 ( .A(instr_jal), .Y(instr_jal_bF_buf0) );
BUFX2 BUFX2_467 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf7_) );
BUFX2 BUFX2_468 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf6_) );
BUFX2 BUFX2_469 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf5_) );
BUFX2 BUFX2_470 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf4_) );
BUFX2 BUFX2_471 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf3_) );
BUFX2 BUFX2_472 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf2_) );
BUFX2 BUFX2_473 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf1_) );
BUFX2 BUFX2_474 ( .A(decoded_rs2_4_), .Y(decoded_rs2_4_bF_buf0_) );
BUFX2 BUFX2_475 ( .A(_5715_), .Y(_5715__bF_buf3) );
BUFX2 BUFX2_476 ( .A(_5715_), .Y(_5715__bF_buf2) );
BUFX2 BUFX2_477 ( .A(_5715_), .Y(_5715__bF_buf1) );
BUFX2 BUFX2_478 ( .A(_5715_), .Y(_5715__bF_buf0) );
BUFX2 BUFX2_479 ( .A(_2173_), .Y(_2173__bF_buf4) );
BUFX2 BUFX2_480 ( .A(_2173_), .Y(_2173__bF_buf3) );
BUFX2 BUFX2_481 ( .A(_2173_), .Y(_2173__bF_buf2) );
BUFX2 BUFX2_482 ( .A(_2173_), .Y(_2173__bF_buf1) );
BUFX2 BUFX2_483 ( .A(_2173_), .Y(_2173__bF_buf0) );
BUFX2 BUFX2_484 ( .A(_4833_), .Y(_4833__bF_buf4) );
BUFX2 BUFX2_485 ( .A(_4833_), .Y(_4833__bF_buf3) );
BUFX2 BUFX2_486 ( .A(_4833_), .Y(_4833__bF_buf2) );
BUFX2 BUFX2_487 ( .A(_4833_), .Y(_4833__bF_buf1) );
BUFX2 BUFX2_488 ( .A(_4833_), .Y(_4833__bF_buf0) );
BUFX2 BUFX2_489 ( .A(_4871_), .Y(_4871__bF_buf4) );
BUFX2 BUFX2_490 ( .A(_4871_), .Y(_4871__bF_buf3) );
BUFX2 BUFX2_491 ( .A(_4871_), .Y(_4871__bF_buf2) );
BUFX2 BUFX2_492 ( .A(_4871_), .Y(_4871__bF_buf1) );
BUFX2 BUFX2_493 ( .A(_4871_), .Y(_4871__bF_buf0) );
BUFX2 BUFX2_494 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf45_) );
BUFX2 BUFX2_495 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf44_) );
BUFX2 BUFX2_496 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf43_) );
BUFX2 BUFX2_497 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf42_) );
BUFX2 BUFX2_498 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf41_) );
BUFX2 BUFX2_499 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf40_) );
BUFX2 BUFX2_500 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf39_) );
BUFX2 BUFX2_501 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf38_) );
BUFX2 BUFX2_502 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf37_) );
BUFX2 BUFX2_503 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf36_) );
BUFX2 BUFX2_504 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf35_) );
BUFX2 BUFX2_505 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf34_) );
BUFX2 BUFX2_506 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf33_) );
BUFX2 BUFX2_507 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf32_) );
BUFX2 BUFX2_508 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf31_) );
BUFX2 BUFX2_509 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf30_) );
BUFX2 BUFX2_510 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf29_) );
BUFX2 BUFX2_511 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf28_) );
BUFX2 BUFX2_512 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf27_) );
BUFX2 BUFX2_513 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf26_) );
BUFX2 BUFX2_514 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf25_) );
BUFX2 BUFX2_515 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf24_) );
BUFX2 BUFX2_516 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf23_) );
BUFX2 BUFX2_517 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf22_) );
BUFX2 BUFX2_518 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf21_) );
BUFX2 BUFX2_519 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf20_) );
BUFX2 BUFX2_520 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf19_) );
BUFX2 BUFX2_521 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf18_) );
BUFX2 BUFX2_522 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf17_) );
BUFX2 BUFX2_523 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf16_) );
BUFX2 BUFX2_524 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf15_) );
BUFX2 BUFX2_525 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf14_) );
BUFX2 BUFX2_526 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf13_) );
BUFX2 BUFX2_527 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf12_) );
BUFX2 BUFX2_528 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf11_) );
BUFX2 BUFX2_529 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf10_) );
BUFX2 BUFX2_530 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf9_) );
BUFX2 BUFX2_531 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf8_) );
BUFX2 BUFX2_532 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf7_) );
BUFX2 BUFX2_533 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf6_) );
BUFX2 BUFX2_534 ( .A(decoded_rs2_1__hier0_bF_buf1), .Y(decoded_rs2_1_bF_buf5_) );
BUFX2 BUFX2_535 ( .A(decoded_rs2_1__hier0_bF_buf0), .Y(decoded_rs2_1_bF_buf4_) );
BUFX2 BUFX2_536 ( .A(decoded_rs2_1__hier0_bF_buf5), .Y(decoded_rs2_1_bF_buf3_) );
BUFX2 BUFX2_537 ( .A(decoded_rs2_1__hier0_bF_buf4), .Y(decoded_rs2_1_bF_buf2_) );
BUFX2 BUFX2_538 ( .A(decoded_rs2_1__hier0_bF_buf3), .Y(decoded_rs2_1_bF_buf1_) );
BUFX2 BUFX2_539 ( .A(decoded_rs2_1__hier0_bF_buf2), .Y(decoded_rs2_1_bF_buf0_) );
BUFX2 BUFX2_540 ( .A(_4639_), .Y(_4639__bF_buf4) );
BUFX2 BUFX2_541 ( .A(_4639_), .Y(_4639__bF_buf3) );
BUFX2 BUFX2_542 ( .A(_4639_), .Y(_4639__bF_buf2) );
BUFX2 BUFX2_543 ( .A(_4639_), .Y(_4639__bF_buf1) );
BUFX2 BUFX2_544 ( .A(_4639_), .Y(_4639__bF_buf0) );
BUFX2 BUFX2_545 ( .A(_7552_), .Y(_7552__bF_buf5) );
BUFX2 BUFX2_546 ( .A(_7552_), .Y(_7552__bF_buf4) );
BUFX2 BUFX2_547 ( .A(_7552_), .Y(_7552__bF_buf3) );
BUFX2 BUFX2_548 ( .A(_7552_), .Y(_7552__bF_buf2) );
BUFX2 BUFX2_549 ( .A(_7552_), .Y(_7552__bF_buf1) );
BUFX2 BUFX2_550 ( .A(_7552_), .Y(_7552__bF_buf0) );
BUFX2 BUFX2_551 ( .A(_4677_), .Y(_4677__bF_buf4) );
BUFX2 BUFX2_552 ( .A(_4677_), .Y(_4677__bF_buf3) );
BUFX2 BUFX2_553 ( .A(_4677_), .Y(_4677__bF_buf2) );
BUFX2 BUFX2_554 ( .A(_4677_), .Y(_4677__bF_buf1) );
BUFX2 BUFX2_555 ( .A(_4677_), .Y(_4677__bF_buf0) );
BUFX2 BUFX2_556 ( .A(_2323_), .Y(_2323__bF_buf3) );
BUFX2 BUFX2_557 ( .A(_2323_), .Y(_2323__bF_buf2) );
BUFX2 BUFX2_558 ( .A(_2323_), .Y(_2323__bF_buf1) );
BUFX2 BUFX2_559 ( .A(_2323_), .Y(_2323__bF_buf0) );
BUFX2 BUFX2_560 ( .A(decoded_rs1_4_), .Y(decoded_rs1_4_bF_buf4_) );
BUFX2 BUFX2_561 ( .A(decoded_rs1_4_), .Y(decoded_rs1_4_bF_buf3_) );
BUFX2 BUFX2_562 ( .A(decoded_rs1_4_), .Y(decoded_rs1_4_bF_buf2_) );
BUFX2 BUFX2_563 ( .A(decoded_rs1_4_), .Y(decoded_rs1_4_bF_buf1_) );
BUFX2 BUFX2_564 ( .A(decoded_rs1_4_), .Y(decoded_rs1_4_bF_buf0_) );
BUFX2 BUFX2_565 ( .A(_2035_), .Y(_2035__bF_buf8) );
BUFX2 BUFX2_566 ( .A(_2035_), .Y(_2035__bF_buf7) );
BUFX2 BUFX2_567 ( .A(_2035_), .Y(_2035__bF_buf6) );
BUFX2 BUFX2_568 ( .A(_2035_), .Y(_2035__bF_buf5) );
BUFX2 BUFX2_569 ( .A(_2035_), .Y(_2035__bF_buf4) );
BUFX2 BUFX2_570 ( .A(_2035_), .Y(_2035__bF_buf3) );
BUFX2 BUFX2_571 ( .A(_2035_), .Y(_2035__bF_buf2) );
BUFX2 BUFX2_572 ( .A(_2035_), .Y(_2035__bF_buf1) );
BUFX2 BUFX2_573 ( .A(_2035_), .Y(_2035__bF_buf0) );
BUFX2 BUFX2_574 ( .A(instr_rdcycle), .Y(instr_rdcycle_bF_buf4) );
BUFX2 BUFX2_575 ( .A(instr_rdcycle), .Y(instr_rdcycle_bF_buf3) );
BUFX2 BUFX2_576 ( .A(instr_rdcycle), .Y(instr_rdcycle_bF_buf2) );
BUFX2 BUFX2_577 ( .A(instr_rdcycle), .Y(instr_rdcycle_bF_buf1) );
BUFX2 BUFX2_578 ( .A(instr_rdcycle), .Y(instr_rdcycle_bF_buf0) );
BUFX2 BUFX2_579 ( .A(_5271_), .Y(_5271__bF_buf3) );
BUFX2 BUFX2_580 ( .A(_5271_), .Y(_5271__bF_buf2) );
BUFX2 BUFX2_581 ( .A(_5271_), .Y(_5271__bF_buf1) );
BUFX2 BUFX2_582 ( .A(_5271_), .Y(_5271__bF_buf0) );
BUFX2 BUFX2_583 ( .A(decoder_pseudo_trigger), .Y(decoder_pseudo_trigger_bF_buf3) );
BUFX2 BUFX2_584 ( .A(decoder_pseudo_trigger), .Y(decoder_pseudo_trigger_bF_buf2) );
BUFX2 BUFX2_585 ( .A(decoder_pseudo_trigger), .Y(decoder_pseudo_trigger_bF_buf1) );
BUFX2 BUFX2_586 ( .A(decoder_pseudo_trigger), .Y(decoder_pseudo_trigger_bF_buf0) );
BUFX2 BUFX2_587 ( .A(_4580_), .Y(_4580__bF_buf4) );
BUFX2 BUFX2_588 ( .A(_4580_), .Y(_4580__bF_buf3) );
BUFX2 BUFX2_589 ( .A(_4580_), .Y(_4580__bF_buf2) );
BUFX2 BUFX2_590 ( .A(_4580_), .Y(_4580__bF_buf1) );
BUFX2 BUFX2_591 ( .A(_4580_), .Y(_4580__bF_buf0) );
BUFX2 BUFX2_592 ( .A(_3011_), .Y(_3011__bF_buf4) );
BUFX2 BUFX2_593 ( .A(_3011_), .Y(_3011__bF_buf3) );
BUFX2 BUFX2_594 ( .A(_3011_), .Y(_3011__bF_buf2) );
BUFX2 BUFX2_595 ( .A(_3011_), .Y(_3011__bF_buf1) );
BUFX2 BUFX2_596 ( .A(_3011_), .Y(_3011__bF_buf0) );
BUFX2 BUFX2_597 ( .A(mem_wordsize_0_), .Y(mem_wordsize_0_bF_buf3_) );
BUFX2 BUFX2_598 ( .A(mem_wordsize_0_), .Y(mem_wordsize_0_bF_buf2_) );
BUFX2 BUFX2_599 ( .A(mem_wordsize_0_), .Y(mem_wordsize_0_bF_buf1_) );
BUFX2 BUFX2_600 ( .A(mem_wordsize_0_), .Y(mem_wordsize_0_bF_buf0_) );
BUFX2 BUFX2_601 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf44_) );
BUFX2 BUFX2_602 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf43_) );
BUFX2 BUFX2_603 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf42_) );
BUFX2 BUFX2_604 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf41_) );
BUFX2 BUFX2_605 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf40_) );
BUFX2 BUFX2_606 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf39_) );
BUFX2 BUFX2_607 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf38_) );
BUFX2 BUFX2_608 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf37_) );
BUFX2 BUFX2_609 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf36_) );
BUFX2 BUFX2_610 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf35_) );
BUFX2 BUFX2_611 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf34_) );
BUFX2 BUFX2_612 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf33_) );
BUFX2 BUFX2_613 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf32_) );
BUFX2 BUFX2_614 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf31_) );
BUFX2 BUFX2_615 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf30_) );
BUFX2 BUFX2_616 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf29_) );
BUFX2 BUFX2_617 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf28_) );
BUFX2 BUFX2_618 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf27_) );
BUFX2 BUFX2_619 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf26_) );
BUFX2 BUFX2_620 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf25_) );
BUFX2 BUFX2_621 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf24_) );
BUFX2 BUFX2_622 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf23_) );
BUFX2 BUFX2_623 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf22_) );
BUFX2 BUFX2_624 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf21_) );
BUFX2 BUFX2_625 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf20_) );
BUFX2 BUFX2_626 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf19_) );
BUFX2 BUFX2_627 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf18_) );
BUFX2 BUFX2_628 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf17_) );
BUFX2 BUFX2_629 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf16_) );
BUFX2 BUFX2_630 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf15_) );
BUFX2 BUFX2_631 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf14_) );
BUFX2 BUFX2_632 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf13_) );
BUFX2 BUFX2_633 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf12_) );
BUFX2 BUFX2_634 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf11_) );
BUFX2 BUFX2_635 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf10_) );
BUFX2 BUFX2_636 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf9_) );
BUFX2 BUFX2_637 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf8_) );
BUFX2 BUFX2_638 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf7_) );
BUFX2 BUFX2_639 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf6_) );
BUFX2 BUFX2_640 ( .A(decoded_rs1_1__hier0_bF_buf2), .Y(decoded_rs1_1_bF_buf5_) );
BUFX2 BUFX2_641 ( .A(decoded_rs1_1__hier0_bF_buf1), .Y(decoded_rs1_1_bF_buf4_) );
BUFX2 BUFX2_642 ( .A(decoded_rs1_1__hier0_bF_buf0), .Y(decoded_rs1_1_bF_buf3_) );
BUFX2 BUFX2_643 ( .A(decoded_rs1_1__hier0_bF_buf5), .Y(decoded_rs1_1_bF_buf2_) );
BUFX2 BUFX2_644 ( .A(decoded_rs1_1__hier0_bF_buf4), .Y(decoded_rs1_1_bF_buf1_) );
BUFX2 BUFX2_645 ( .A(decoded_rs1_1__hier0_bF_buf3), .Y(decoded_rs1_1_bF_buf0_) );
BUFX2 BUFX2_646 ( .A(_4539_), .Y(_4539__bF_buf3) );
BUFX2 BUFX2_647 ( .A(_4539_), .Y(_4539__bF_buf2) );
BUFX2 BUFX2_648 ( .A(_4539_), .Y(_4539__bF_buf1) );
BUFX2 BUFX2_649 ( .A(_4539_), .Y(_4539__bF_buf0) );
BUFX2 BUFX2_650 ( .A(_1817_), .Y(_1817__bF_buf3) );
BUFX2 BUFX2_651 ( .A(_1817_), .Y(_1817__bF_buf2) );
BUFX2 BUFX2_652 ( .A(_1817_), .Y(_1817__bF_buf1) );
BUFX2 BUFX2_653 ( .A(_1817_), .Y(_1817__bF_buf0) );
BUFX2 BUFX2_654 ( .A(_5706_), .Y(_5706__bF_buf11) );
BUFX2 BUFX2_655 ( .A(_5706_), .Y(_5706__bF_buf10) );
BUFX2 BUFX2_656 ( .A(_5706_), .Y(_5706__bF_buf9) );
BUFX2 BUFX2_657 ( .A(_5706_), .Y(_5706__bF_buf8) );
BUFX2 BUFX2_658 ( .A(_5706_), .Y(_5706__bF_buf7) );
BUFX2 BUFX2_659 ( .A(_5706_), .Y(_5706__bF_buf6) );
BUFX2 BUFX2_660 ( .A(_5706_), .Y(_5706__bF_buf5) );
BUFX2 BUFX2_661 ( .A(_5706_), .Y(_5706__bF_buf4) );
BUFX2 BUFX2_662 ( .A(_5706_), .Y(_5706__bF_buf3) );
BUFX2 BUFX2_663 ( .A(_5706_), .Y(_5706__bF_buf2) );
BUFX2 BUFX2_664 ( .A(_5706_), .Y(_5706__bF_buf1) );
BUFX2 BUFX2_665 ( .A(_5706_), .Y(_5706__bF_buf0) );
BUFX2 BUFX2_666 ( .A(_3810_), .Y(_3810__bF_buf4) );
BUFX2 BUFX2_667 ( .A(_3810_), .Y(_3810__bF_buf3) );
BUFX2 BUFX2_668 ( .A(_3810_), .Y(_3810__bF_buf2) );
BUFX2 BUFX2_669 ( .A(_3810_), .Y(_3810__bF_buf1) );
BUFX2 BUFX2_670 ( .A(_3810_), .Y(_3810__bF_buf0) );
BUFX2 BUFX2_671 ( .A(_4824_), .Y(_4824__bF_buf4) );
BUFX2 BUFX2_672 ( .A(_4824_), .Y(_4824__bF_buf3) );
BUFX2 BUFX2_673 ( .A(_4824_), .Y(_4824__bF_buf2) );
BUFX2 BUFX2_674 ( .A(_4824_), .Y(_4824__bF_buf1) );
BUFX2 BUFX2_675 ( .A(_4824_), .Y(_4824__bF_buf0) );
BUFX2 BUFX2_676 ( .A(_5362_), .Y(_5362__bF_buf14) );
BUFX2 BUFX2_677 ( .A(_5362_), .Y(_5362__bF_buf13) );
BUFX2 BUFX2_678 ( .A(_5362_), .Y(_5362__bF_buf12) );
BUFX2 BUFX2_679 ( .A(_5362_), .Y(_5362__bF_buf11) );
BUFX2 BUFX2_680 ( .A(_5362_), .Y(_5362__bF_buf10) );
BUFX2 BUFX2_681 ( .A(_5362_), .Y(_5362__bF_buf9) );
BUFX2 BUFX2_682 ( .A(_5362_), .Y(_5362__bF_buf8) );
BUFX2 BUFX2_683 ( .A(_5362_), .Y(_5362__bF_buf7) );
BUFX2 BUFX2_684 ( .A(_5362_), .Y(_5362__bF_buf6) );
BUFX2 BUFX2_685 ( .A(_5362_), .Y(_5362__bF_buf5) );
BUFX2 BUFX2_686 ( .A(_5362_), .Y(_5362__bF_buf4) );
BUFX2 BUFX2_687 ( .A(_5362_), .Y(_5362__bF_buf3) );
BUFX2 BUFX2_688 ( .A(_5362_), .Y(_5362__bF_buf2) );
BUFX2 BUFX2_689 ( .A(_5362_), .Y(_5362__bF_buf1) );
BUFX2 BUFX2_690 ( .A(_5362_), .Y(_5362__bF_buf0) );
BUFX2 BUFX2_691 ( .A(_10728__2_), .Y(_10728__2_bF_buf4_) );
BUFX2 BUFX2_692 ( .A(_10728__2_), .Y(_10728__2_bF_buf3_) );
BUFX2 BUFX2_693 ( .A(_10728__2_), .Y(_10728__2_bF_buf2_) );
BUFX2 BUFX2_694 ( .A(_10728__2_), .Y(_10728__2_bF_buf1_) );
BUFX2 BUFX2_695 ( .A(_10728__2_), .Y(_10728__2_bF_buf0_) );
BUFX2 BUFX2_696 ( .A(_3005_), .Y(_3005__bF_buf4) );
BUFX2 BUFX2_697 ( .A(_3005_), .Y(_3005__bF_buf3) );
BUFX2 BUFX2_698 ( .A(_3005_), .Y(_3005__bF_buf2) );
BUFX2 BUFX2_699 ( .A(_3005_), .Y(_3005__bF_buf1) );
BUFX2 BUFX2_700 ( .A(_3005_), .Y(_3005__bF_buf0) );
BUFX2 BUFX2_701 ( .A(_4439_), .Y(_4439__bF_buf6) );
BUFX2 BUFX2_702 ( .A(_4439_), .Y(_4439__bF_buf5) );
BUFX2 BUFX2_703 ( .A(_4439_), .Y(_4439__bF_buf4) );
BUFX2 BUFX2_704 ( .A(_4439_), .Y(_4439__bF_buf3) );
BUFX2 BUFX2_705 ( .A(_4439_), .Y(_4439__bF_buf2) );
BUFX2 BUFX2_706 ( .A(_4439_), .Y(_4439__bF_buf1) );
BUFX2 BUFX2_707 ( .A(_4439_), .Y(_4439__bF_buf0) );
BUFX2 BUFX2_708 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf5_) );
BUFX2 BUFX2_709 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf4_) );
BUFX2 BUFX2_710 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf3_) );
BUFX2 BUFX2_711 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf2_) );
BUFX2 BUFX2_712 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf1_) );
BUFX2 BUFX2_713 ( .A(cpu_state_1_), .Y(cpu_state_1_bF_buf0_) );
BUFX2 BUFX2_714 ( .A(_3880_), .Y(_3880__bF_buf7) );
BUFX2 BUFX2_715 ( .A(_3880_), .Y(_3880__bF_buf6) );
BUFX2 BUFX2_716 ( .A(_3880_), .Y(_3880__bF_buf5) );
BUFX2 BUFX2_717 ( .A(_3880_), .Y(_3880__bF_buf4) );
BUFX2 BUFX2_718 ( .A(_3880_), .Y(_3880__bF_buf3) );
BUFX2 BUFX2_719 ( .A(_3880_), .Y(_3880__bF_buf2) );
BUFX2 BUFX2_720 ( .A(_3880_), .Y(_3880__bF_buf1) );
BUFX2 BUFX2_721 ( .A(_3880_), .Y(_3880__bF_buf0) );
BUFX2 BUFX2_722 ( .A(_7631_), .Y(_7631__bF_buf5) );
BUFX2 BUFX2_723 ( .A(_7631_), .Y(_7631__bF_buf4) );
BUFX2 BUFX2_724 ( .A(_7631_), .Y(_7631__bF_buf3) );
BUFX2 BUFX2_725 ( .A(_7631_), .Y(_7631__bF_buf2) );
BUFX2 BUFX2_726 ( .A(_7631_), .Y(_7631__bF_buf1) );
BUFX2 BUFX2_727 ( .A(_7631_), .Y(_7631__bF_buf0) );
BUFX2 BUFX2_728 ( .A(_4985_), .Y(_4985__bF_buf8) );
BUFX2 BUFX2_729 ( .A(_4985_), .Y(_4985__bF_buf7) );
BUFX2 BUFX2_730 ( .A(_4985_), .Y(_4985__bF_buf6) );
BUFX2 BUFX2_731 ( .A(_4985_), .Y(_4985__bF_buf5) );
BUFX2 BUFX2_732 ( .A(_4985_), .Y(_4985__bF_buf4) );
BUFX2 BUFX2_733 ( .A(_4985_), .Y(_4985__bF_buf3) );
BUFX2 BUFX2_734 ( .A(_4985_), .Y(_4985__bF_buf2) );
BUFX2 BUFX2_735 ( .A(_4985_), .Y(_4985__bF_buf1) );
BUFX2 BUFX2_736 ( .A(_4985_), .Y(_4985__bF_buf0) );
BUFX2 BUFX2_737 ( .A(_4621_), .Y(_4621__bF_buf4) );
BUFX2 BUFX2_738 ( .A(_4621_), .Y(_4621__bF_buf3) );
BUFX2 BUFX2_739 ( .A(_4621_), .Y(_4621__bF_buf2) );
BUFX2 BUFX2_740 ( .A(_4621_), .Y(_4621__bF_buf1) );
BUFX2 BUFX2_741 ( .A(_4621_), .Y(_4621__bF_buf0) );
BUFX2 BUFX2_742 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf48) );
BUFX2 BUFX2_743 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf47) );
BUFX2 BUFX2_744 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf46) );
BUFX2 BUFX2_745 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf45) );
BUFX2 BUFX2_746 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf44) );
BUFX2 BUFX2_747 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf43) );
BUFX2 BUFX2_748 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf42) );
BUFX2 BUFX2_749 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf41) );
BUFX2 BUFX2_750 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf40) );
BUFX2 BUFX2_751 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf39) );
BUFX2 BUFX2_752 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf38) );
BUFX2 BUFX2_753 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf37) );
BUFX2 BUFX2_754 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf36) );
BUFX2 BUFX2_755 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf35) );
BUFX2 BUFX2_756 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf34) );
BUFX2 BUFX2_757 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf33) );
BUFX2 BUFX2_758 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf32) );
BUFX2 BUFX2_759 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf31) );
BUFX2 BUFX2_760 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf30) );
BUFX2 BUFX2_761 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf29) );
BUFX2 BUFX2_762 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf28) );
BUFX2 BUFX2_763 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf27) );
BUFX2 BUFX2_764 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf26) );
BUFX2 BUFX2_765 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf25) );
BUFX2 BUFX2_766 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf24) );
BUFX2 BUFX2_767 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf23) );
BUFX2 BUFX2_768 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf22) );
BUFX2 BUFX2_769 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf21) );
BUFX2 BUFX2_770 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf20) );
BUFX2 BUFX2_771 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf19) );
BUFX2 BUFX2_772 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf18) );
BUFX2 BUFX2_773 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf17) );
BUFX2 BUFX2_774 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf16) );
BUFX2 BUFX2_775 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf15) );
BUFX2 BUFX2_776 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf14) );
BUFX2 BUFX2_777 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf13) );
BUFX2 BUFX2_778 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf12) );
BUFX2 BUFX2_779 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf11) );
BUFX2 BUFX2_780 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf10) );
BUFX2 BUFX2_781 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf9) );
BUFX2 BUFX2_782 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf8) );
BUFX2 BUFX2_783 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf7) );
BUFX2 BUFX2_784 ( .A(_7569__hier0_bF_buf6), .Y(_7569__bF_buf6) );
BUFX2 BUFX2_785 ( .A(_7569__hier0_bF_buf5), .Y(_7569__bF_buf5) );
BUFX2 BUFX2_786 ( .A(_7569__hier0_bF_buf4), .Y(_7569__bF_buf4) );
BUFX2 BUFX2_787 ( .A(_7569__hier0_bF_buf3), .Y(_7569__bF_buf3) );
BUFX2 BUFX2_788 ( .A(_7569__hier0_bF_buf2), .Y(_7569__bF_buf2) );
BUFX2 BUFX2_789 ( .A(_7569__hier0_bF_buf1), .Y(_7569__bF_buf1) );
BUFX2 BUFX2_790 ( .A(_7569__hier0_bF_buf0), .Y(_7569__bF_buf0) );
BUFX2 BUFX2_791 ( .A(_2378_), .Y(_2378__bF_buf7) );
BUFX2 BUFX2_792 ( .A(_2378_), .Y(_2378__bF_buf6) );
BUFX2 BUFX2_793 ( .A(_2378_), .Y(_2378__bF_buf5) );
BUFX2 BUFX2_794 ( .A(_2378_), .Y(_2378__bF_buf4) );
BUFX2 BUFX2_795 ( .A(_2378_), .Y(_2378__bF_buf3) );
BUFX2 BUFX2_796 ( .A(_2378_), .Y(_2378__bF_buf2) );
BUFX2 BUFX2_797 ( .A(_2378_), .Y(_2378__bF_buf1) );
BUFX2 BUFX2_798 ( .A(_2378_), .Y(_2378__bF_buf0) );
BUFX2 BUFX2_799 ( .A(instr_rdcycleh), .Y(instr_rdcycleh_bF_buf3) );
BUFX2 BUFX2_800 ( .A(instr_rdcycleh), .Y(instr_rdcycleh_bF_buf2) );
BUFX2 BUFX2_801 ( .A(instr_rdcycleh), .Y(instr_rdcycleh_bF_buf1) );
BUFX2 BUFX2_802 ( .A(instr_rdcycleh), .Y(instr_rdcycleh_bF_buf0) );
BUFX2 BUFX2_803 ( .A(_4597_), .Y(_4597__bF_buf3) );
BUFX2 BUFX2_804 ( .A(_4597_), .Y(_4597__bF_buf2) );
BUFX2 BUFX2_805 ( .A(_4597_), .Y(_4597__bF_buf1) );
BUFX2 BUFX2_806 ( .A(_4597_), .Y(_4597__bF_buf0) );
BUFX2 BUFX2_807 ( .A(_4806_), .Y(_4806__bF_buf4) );
BUFX2 BUFX2_808 ( .A(_4806_), .Y(_4806__bF_buf3) );
BUFX2 BUFX2_809 ( .A(_4806_), .Y(_4806__bF_buf2) );
BUFX2 BUFX2_810 ( .A(_4806_), .Y(_4806__bF_buf1) );
BUFX2 BUFX2_811 ( .A(_4806_), .Y(_4806__bF_buf0) );
BUFX2 BUFX2_812 ( .A(_7698_), .Y(_7698__bF_buf4) );
BUFX2 BUFX2_813 ( .A(_7698_), .Y(_7698__bF_buf3) );
BUFX2 BUFX2_814 ( .A(_7698_), .Y(_7698__bF_buf2) );
BUFX2 BUFX2_815 ( .A(_7698_), .Y(_7698__bF_buf1) );
BUFX2 BUFX2_816 ( .A(_7698_), .Y(_7698__bF_buf0) );
BUFX2 BUFX2_817 ( .A(_4747_), .Y(_4747__bF_buf4) );
BUFX2 BUFX2_818 ( .A(_4747_), .Y(_4747__bF_buf3) );
BUFX2 BUFX2_819 ( .A(_4747_), .Y(_4747__bF_buf2) );
BUFX2 BUFX2_820 ( .A(_4747_), .Y(_4747__bF_buf1) );
BUFX2 BUFX2_821 ( .A(_4747_), .Y(_4747__bF_buf0) );
BUFX2 BUFX2_822 ( .A(_4080_), .Y(_4080__bF_buf7) );
BUFX2 BUFX2_823 ( .A(_4080_), .Y(_4080__bF_buf6) );
BUFX2 BUFX2_824 ( .A(_4080_), .Y(_4080__bF_buf5) );
BUFX2 BUFX2_825 ( .A(_4080_), .Y(_4080__bF_buf4) );
BUFX2 BUFX2_826 ( .A(_4080_), .Y(_4080__bF_buf3) );
BUFX2 BUFX2_827 ( .A(_4080_), .Y(_4080__bF_buf2) );
BUFX2 BUFX2_828 ( .A(_4080_), .Y(_4080__bF_buf1) );
BUFX2 BUFX2_829 ( .A(_4080_), .Y(_4080__bF_buf0) );
BUFX2 BUFX2_830 ( .A(_2240_), .Y(_2240__bF_buf7) );
BUFX2 BUFX2_831 ( .A(_2240_), .Y(_2240__bF_buf6) );
BUFX2 BUFX2_832 ( .A(_2240_), .Y(_2240__bF_buf5) );
BUFX2 BUFX2_833 ( .A(_2240_), .Y(_2240__bF_buf4) );
BUFX2 BUFX2_834 ( .A(_2240_), .Y(_2240__bF_buf3) );
BUFX2 BUFX2_835 ( .A(_2240_), .Y(_2240__bF_buf2) );
BUFX2 BUFX2_836 ( .A(_2240_), .Y(_2240__bF_buf1) );
BUFX2 BUFX2_837 ( .A(_2240_), .Y(_2240__bF_buf0) );
BUFX2 BUFX2_838 ( .A(resetn), .Y(resetn_bF_buf11) );
BUFX2 BUFX2_839 ( .A(resetn), .Y(resetn_bF_buf10) );
BUFX2 BUFX2_840 ( .A(resetn), .Y(resetn_bF_buf9) );
BUFX2 BUFX2_841 ( .A(resetn), .Y(resetn_bF_buf8) );
BUFX2 BUFX2_842 ( .A(resetn), .Y(resetn_bF_buf7) );
BUFX2 BUFX2_843 ( .A(resetn), .Y(resetn_bF_buf6) );
BUFX2 BUFX2_844 ( .A(resetn), .Y(resetn_bF_buf5) );
BUFX2 BUFX2_845 ( .A(resetn), .Y(resetn_bF_buf4) );
BUFX2 BUFX2_846 ( .A(resetn), .Y(resetn_bF_buf3) );
BUFX2 BUFX2_847 ( .A(resetn), .Y(resetn_bF_buf2) );
BUFX2 BUFX2_848 ( .A(resetn), .Y(resetn_bF_buf1) );
BUFX2 BUFX2_849 ( .A(resetn), .Y(resetn_bF_buf0) );
BUFX2 BUFX2_850 ( .A(_7560_), .Y(_7560__bF_buf12) );
BUFX2 BUFX2_851 ( .A(_7560_), .Y(_7560__bF_buf11) );
BUFX2 BUFX2_852 ( .A(_7560_), .Y(_7560__bF_buf10) );
BUFX2 BUFX2_853 ( .A(_7560_), .Y(_7560__bF_buf9) );
BUFX2 BUFX2_854 ( .A(_7560_), .Y(_7560__bF_buf8) );
BUFX2 BUFX2_855 ( .A(_7560_), .Y(_7560__bF_buf7) );
BUFX2 BUFX2_856 ( .A(_7560_), .Y(_7560__bF_buf6) );
BUFX2 BUFX2_857 ( .A(_7560_), .Y(_7560__bF_buf5) );
BUFX2 BUFX2_858 ( .A(_7560_), .Y(_7560__bF_buf4) );
BUFX2 BUFX2_859 ( .A(_7560_), .Y(_7560__bF_buf3) );
BUFX2 BUFX2_860 ( .A(_7560_), .Y(_7560__bF_buf2) );
BUFX2 BUFX2_861 ( .A(_7560_), .Y(_7560__bF_buf1) );
BUFX2 BUFX2_862 ( .A(_7560_), .Y(_7560__bF_buf0) );
BUFX2 BUFX2_863 ( .A(_4685_), .Y(_4685__bF_buf4) );
BUFX2 BUFX2_864 ( .A(_4685_), .Y(_4685__bF_buf3) );
BUFX2 BUFX2_865 ( .A(_4685_), .Y(_4685__bF_buf2) );
BUFX2 BUFX2_866 ( .A(_4685_), .Y(_4685__bF_buf1) );
BUFX2 BUFX2_867 ( .A(_4685_), .Y(_4685__bF_buf0) );
BUFX2 BUFX2_868 ( .A(_4703_), .Y(_4703__bF_buf4) );
BUFX2 BUFX2_869 ( .A(_4703_), .Y(_4703__bF_buf3) );
BUFX2 BUFX2_870 ( .A(_4703_), .Y(_4703__bF_buf2) );
BUFX2 BUFX2_871 ( .A(_4703_), .Y(_4703__bF_buf1) );
BUFX2 BUFX2_872 ( .A(_4703_), .Y(_4703__bF_buf0) );
BUFX2 BUFX2_873 ( .A(_5890_), .Y(_5890__bF_buf3) );
BUFX2 BUFX2_874 ( .A(_5890_), .Y(_5890__bF_buf2) );
BUFX2 BUFX2_875 ( .A(_5890_), .Y(_5890__bF_buf1) );
BUFX2 BUFX2_876 ( .A(_5890_), .Y(_5890__bF_buf0) );
BUFX2 BUFX2_877 ( .A(_10118_), .Y(_10118__bF_buf4) );
BUFX2 BUFX2_878 ( .A(_10118_), .Y(_10118__bF_buf3) );
BUFX2 BUFX2_879 ( .A(_10118_), .Y(_10118__bF_buf2) );
BUFX2 BUFX2_880 ( .A(_10118_), .Y(_10118__bF_buf1) );
BUFX2 BUFX2_881 ( .A(_10118_), .Y(_10118__bF_buf0) );
BUFX2 BUFX2_882 ( .A(instr_sub), .Y(instr_sub_bF_buf4) );
BUFX2 BUFX2_883 ( .A(instr_sub), .Y(instr_sub_bF_buf3) );
BUFX2 BUFX2_884 ( .A(instr_sub), .Y(instr_sub_bF_buf2) );
BUFX2 BUFX2_885 ( .A(instr_sub), .Y(instr_sub_bF_buf1) );
BUFX2 BUFX2_886 ( .A(instr_sub), .Y(instr_sub_bF_buf0) );
BUFX2 BUFX2_887 ( .A(_5849_), .Y(_5849__bF_buf4) );
BUFX2 BUFX2_888 ( .A(_5849_), .Y(_5849__bF_buf3) );
BUFX2 BUFX2_889 ( .A(_5849_), .Y(_5849__bF_buf2) );
BUFX2 BUFX2_890 ( .A(_5849_), .Y(_5849__bF_buf1) );
BUFX2 BUFX2_891 ( .A(_5849_), .Y(_5849__bF_buf0) );
BUFX2 BUFX2_892 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf5) );
BUFX2 BUFX2_893 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf4) );
BUFX2 BUFX2_894 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf3) );
BUFX2 BUFX2_895 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf2) );
BUFX2 BUFX2_896 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf1) );
BUFX2 BUFX2_897 ( .A(mem_do_prefetch), .Y(mem_do_prefetch_bF_buf0) );
BUFX2 BUFX2_898 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf6_) );
BUFX2 BUFX2_899 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf5_) );
BUFX2 BUFX2_900 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf4_) );
BUFX2 BUFX2_901 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf3_) );
BUFX2 BUFX2_902 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf2_) );
BUFX2 BUFX2_903 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf1_) );
BUFX2 BUFX2_904 ( .A(decoded_rs2_3_), .Y(decoded_rs2_3_bF_buf0_) );
BUFX2 BUFX2_905 ( .A(_2037_), .Y(_2037__bF_buf4) );
BUFX2 BUFX2_906 ( .A(_2037_), .Y(_2037__bF_buf3) );
BUFX2 BUFX2_907 ( .A(_2037_), .Y(_2037__bF_buf2) );
BUFX2 BUFX2_908 ( .A(_2037_), .Y(_2037__bF_buf1) );
BUFX2 BUFX2_909 ( .A(_2037_), .Y(_2037__bF_buf0) );
BUFX2 BUFX2_910 ( .A(mem_do_rinst), .Y(mem_do_rinst_bF_buf4) );
BUFX2 BUFX2_911 ( .A(mem_do_rinst), .Y(mem_do_rinst_bF_buf3) );
BUFX2 BUFX2_912 ( .A(mem_do_rinst), .Y(mem_do_rinst_bF_buf2) );
BUFX2 BUFX2_913 ( .A(mem_do_rinst), .Y(mem_do_rinst_bF_buf1) );
BUFX2 BUFX2_914 ( .A(mem_do_rinst), .Y(mem_do_rinst_bF_buf0) );
BUFX2 BUFX2_915 ( .A(_4641_), .Y(_4641__bF_buf6) );
BUFX2 BUFX2_916 ( .A(_4641_), .Y(_4641__bF_buf5) );
BUFX2 BUFX2_917 ( .A(_4641_), .Y(_4641__bF_buf4) );
BUFX2 BUFX2_918 ( .A(_4641_), .Y(_4641__bF_buf3) );
BUFX2 BUFX2_919 ( .A(_4641_), .Y(_4641__bF_buf2) );
BUFX2 BUFX2_920 ( .A(_4641_), .Y(_4641__bF_buf1) );
BUFX2 BUFX2_921 ( .A(_4641_), .Y(_4641__bF_buf0) );
BUFX2 BUFX2_922 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf78_) );
BUFX2 BUFX2_923 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf77_) );
BUFX2 BUFX2_924 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf76_) );
BUFX2 BUFX2_925 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf75_) );
BUFX2 BUFX2_926 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf74_) );
BUFX2 BUFX2_927 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf73_) );
BUFX2 BUFX2_928 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf72_) );
BUFX2 BUFX2_929 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf71_) );
BUFX2 BUFX2_930 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf70_) );
BUFX2 BUFX2_931 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf69_) );
BUFX2 BUFX2_932 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf68_) );
BUFX2 BUFX2_933 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf67_) );
BUFX2 BUFX2_934 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf66_) );
BUFX2 BUFX2_935 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf65_) );
BUFX2 BUFX2_936 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf64_) );
BUFX2 BUFX2_937 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf63_) );
BUFX2 BUFX2_938 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf62_) );
BUFX2 BUFX2_939 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf61_) );
BUFX2 BUFX2_940 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf60_) );
BUFX2 BUFX2_941 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf59_) );
BUFX2 BUFX2_942 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf58_) );
BUFX2 BUFX2_943 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf57_) );
BUFX2 BUFX2_944 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf56_) );
BUFX2 BUFX2_945 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf55_) );
BUFX2 BUFX2_946 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf54_) );
BUFX2 BUFX2_947 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf53_) );
BUFX2 BUFX2_948 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf52_) );
BUFX2 BUFX2_949 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf51_) );
BUFX2 BUFX2_950 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf50_) );
BUFX2 BUFX2_951 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf49_) );
BUFX2 BUFX2_952 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf48_) );
BUFX2 BUFX2_953 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf47_) );
BUFX2 BUFX2_954 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf46_) );
BUFX2 BUFX2_955 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf45_) );
BUFX2 BUFX2_956 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf44_) );
BUFX2 BUFX2_957 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf43_) );
BUFX2 BUFX2_958 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf42_) );
BUFX2 BUFX2_959 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf41_) );
BUFX2 BUFX2_960 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf40_) );
BUFX2 BUFX2_961 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf39_) );
BUFX2 BUFX2_962 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf38_) );
BUFX2 BUFX2_963 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf37_) );
BUFX2 BUFX2_964 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf36_) );
BUFX2 BUFX2_965 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf35_) );
BUFX2 BUFX2_966 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf34_) );
BUFX2 BUFX2_967 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf33_) );
BUFX2 BUFX2_968 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf32_) );
BUFX2 BUFX2_969 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf31_) );
BUFX2 BUFX2_970 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf30_) );
BUFX2 BUFX2_971 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf29_) );
BUFX2 BUFX2_972 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf28_) );
BUFX2 BUFX2_973 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf27_) );
BUFX2 BUFX2_974 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf26_) );
BUFX2 BUFX2_975 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf25_) );
BUFX2 BUFX2_976 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf24_) );
BUFX2 BUFX2_977 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf23_) );
BUFX2 BUFX2_978 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf22_) );
BUFX2 BUFX2_979 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf21_) );
BUFX2 BUFX2_980 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf20_) );
BUFX2 BUFX2_981 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf19_) );
BUFX2 BUFX2_982 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf18_) );
BUFX2 BUFX2_983 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf17_) );
BUFX2 BUFX2_984 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf16_) );
BUFX2 BUFX2_985 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf15_) );
BUFX2 BUFX2_986 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf14_) );
BUFX2 BUFX2_987 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf13_) );
BUFX2 BUFX2_988 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf12_) );
BUFX2 BUFX2_989 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf11_) );
BUFX2 BUFX2_990 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf10_) );
BUFX2 BUFX2_991 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf9_) );
BUFX2 BUFX2_992 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf8_) );
BUFX2 BUFX2_993 ( .A(decoded_rs2_0__hier0_bF_buf0), .Y(decoded_rs2_0_bF_buf7_) );
BUFX2 BUFX2_994 ( .A(decoded_rs2_0__hier0_bF_buf7), .Y(decoded_rs2_0_bF_buf6_) );
BUFX2 BUFX2_995 ( .A(decoded_rs2_0__hier0_bF_buf6), .Y(decoded_rs2_0_bF_buf5_) );
BUFX2 BUFX2_996 ( .A(decoded_rs2_0__hier0_bF_buf5), .Y(decoded_rs2_0_bF_buf4_) );
BUFX2 BUFX2_997 ( .A(decoded_rs2_0__hier0_bF_buf4), .Y(decoded_rs2_0_bF_buf3_) );
BUFX2 BUFX2_998 ( .A(decoded_rs2_0__hier0_bF_buf3), .Y(decoded_rs2_0_bF_buf2_) );
BUFX2 BUFX2_999 ( .A(decoded_rs2_0__hier0_bF_buf2), .Y(decoded_rs2_0_bF_buf1_) );
BUFX2 BUFX2_1000 ( .A(decoded_rs2_0__hier0_bF_buf1), .Y(decoded_rs2_0_bF_buf0_) );
BUFX2 BUFX2_1001 ( .A(_4447_), .Y(_4447__bF_buf3) );
BUFX2 BUFX2_1002 ( .A(_4447_), .Y(_4447__bF_buf2) );
BUFX2 BUFX2_1003 ( .A(_4447_), .Y(_4447__bF_buf1) );
BUFX2 BUFX2_1004 ( .A(_4447_), .Y(_4447__bF_buf0) );
BUFX2 BUFX2_1005 ( .A(_7551_), .Y(_7551__bF_buf3) );
BUFX2 BUFX2_1006 ( .A(_7551_), .Y(_7551__bF_buf2) );
BUFX2 BUFX2_1007 ( .A(_7551_), .Y(_7551__bF_buf1) );
BUFX2 BUFX2_1008 ( .A(_7551_), .Y(_7551__bF_buf0) );
BUFX2 BUFX2_1009 ( .A(_3947_), .Y(_3947__bF_buf7) );
BUFX2 BUFX2_1010 ( .A(_3947_), .Y(_3947__bF_buf6) );
BUFX2 BUFX2_1011 ( .A(_3947_), .Y(_3947__bF_buf5) );
BUFX2 BUFX2_1012 ( .A(_3947_), .Y(_3947__bF_buf4) );
BUFX2 BUFX2_1013 ( .A(_3947_), .Y(_3947__bF_buf3) );
BUFX2 BUFX2_1014 ( .A(_3947_), .Y(_3947__bF_buf2) );
BUFX2 BUFX2_1015 ( .A(_3947_), .Y(_3947__bF_buf1) );
BUFX2 BUFX2_1016 ( .A(_3947_), .Y(_3947__bF_buf0) );
BUFX2 BUFX2_1017 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf6_) );
BUFX2 BUFX2_1018 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf5_) );
BUFX2 BUFX2_1019 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf4_) );
BUFX2 BUFX2_1020 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf3_) );
BUFX2 BUFX2_1021 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf2_) );
BUFX2 BUFX2_1022 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf1_) );
BUFX2 BUFX2_1023 ( .A(decoded_rs1_3_), .Y(decoded_rs1_3_bF_buf0_) );
BUFX2 BUFX2_1024 ( .A(_4579_), .Y(_4579__bF_buf4) );
BUFX2 BUFX2_1025 ( .A(_4579_), .Y(_4579__bF_buf3) );
BUFX2 BUFX2_1026 ( .A(_4579_), .Y(_4579__bF_buf2) );
BUFX2 BUFX2_1027 ( .A(_4579_), .Y(_4579__bF_buf1) );
BUFX2 BUFX2_1028 ( .A(_4579_), .Y(_4579__bF_buf0) );
BUFX2 BUFX2_1029 ( .A(_7586_), .Y(_7586__bF_buf3) );
BUFX2 BUFX2_1030 ( .A(_7586_), .Y(_7586__bF_buf2) );
BUFX2 BUFX2_1031 ( .A(_7586_), .Y(_7586__bF_buf1) );
BUFX2 BUFX2_1032 ( .A(_7586_), .Y(_7586__bF_buf0) );
BUFX2 BUFX2_1033 ( .A(_5746_), .Y(_5746__bF_buf7) );
BUFX2 BUFX2_1034 ( .A(_5746_), .Y(_5746__bF_buf6) );
BUFX2 BUFX2_1035 ( .A(_5746_), .Y(_5746__bF_buf5) );
BUFX2 BUFX2_1036 ( .A(_5746_), .Y(_5746__bF_buf4) );
BUFX2 BUFX2_1037 ( .A(_5746_), .Y(_5746__bF_buf3) );
BUFX2 BUFX2_1038 ( .A(_5746_), .Y(_5746__bF_buf2) );
BUFX2 BUFX2_1039 ( .A(_5746_), .Y(_5746__bF_buf1) );
BUFX2 BUFX2_1040 ( .A(_5746_), .Y(_5746__bF_buf0) );
BUFX2 BUFX2_1041 ( .A(_10109_), .Y(_10109__bF_buf4) );
BUFX2 BUFX2_1042 ( .A(_10109_), .Y(_10109__bF_buf3) );
BUFX2 BUFX2_1043 ( .A(_10109_), .Y(_10109__bF_buf2) );
BUFX2 BUFX2_1044 ( .A(_10109_), .Y(_10109__bF_buf1) );
BUFX2 BUFX2_1045 ( .A(_10109_), .Y(_10109__bF_buf0) );
BUFX2 BUFX2_1046 ( .A(_10728__4_), .Y(_10728__4_bF_buf4_) );
BUFX2 BUFX2_1047 ( .A(_10728__4_), .Y(_10728__4_bF_buf3_) );
BUFX2 BUFX2_1048 ( .A(_10728__4_), .Y(_10728__4_bF_buf2_) );
BUFX2 BUFX2_1049 ( .A(_10728__4_), .Y(_10728__4_bF_buf1_) );
BUFX2 BUFX2_1050 ( .A(_10728__4_), .Y(_10728__4_bF_buf0_) );
BUFX2 BUFX2_1051 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf57_) );
BUFX2 BUFX2_1052 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf56_) );
BUFX2 BUFX2_1053 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf55_) );
BUFX2 BUFX2_1054 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf54_) );
BUFX2 BUFX2_1055 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf53_) );
BUFX2 BUFX2_1056 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf52_) );
BUFX2 BUFX2_1057 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf51_) );
BUFX2 BUFX2_1058 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf50_) );
BUFX2 BUFX2_1059 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf49_) );
BUFX2 BUFX2_1060 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf48_) );
BUFX2 BUFX2_1061 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf47_) );
BUFX2 BUFX2_1062 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf46_) );
BUFX2 BUFX2_1063 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf45_) );
BUFX2 BUFX2_1064 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf44_) );
BUFX2 BUFX2_1065 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf43_) );
BUFX2 BUFX2_1066 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf42_) );
BUFX2 BUFX2_1067 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf41_) );
BUFX2 BUFX2_1068 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf40_) );
BUFX2 BUFX2_1069 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf39_) );
BUFX2 BUFX2_1070 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf38_) );
BUFX2 BUFX2_1071 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf37_) );
BUFX2 BUFX2_1072 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf36_) );
BUFX2 BUFX2_1073 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf35_) );
BUFX2 BUFX2_1074 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf34_) );
BUFX2 BUFX2_1075 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf33_) );
BUFX2 BUFX2_1076 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf32_) );
BUFX2 BUFX2_1077 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf31_) );
BUFX2 BUFX2_1078 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf30_) );
BUFX2 BUFX2_1079 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf29_) );
BUFX2 BUFX2_1080 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf28_) );
BUFX2 BUFX2_1081 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf27_) );
BUFX2 BUFX2_1082 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf26_) );
BUFX2 BUFX2_1083 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf25_) );
BUFX2 BUFX2_1084 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf24_) );
BUFX2 BUFX2_1085 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf23_) );
BUFX2 BUFX2_1086 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf22_) );
BUFX2 BUFX2_1087 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf21_) );
BUFX2 BUFX2_1088 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf20_) );
BUFX2 BUFX2_1089 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf19_) );
BUFX2 BUFX2_1090 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf18_) );
BUFX2 BUFX2_1091 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf17_) );
BUFX2 BUFX2_1092 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf16_) );
BUFX2 BUFX2_1093 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf15_) );
BUFX2 BUFX2_1094 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf14_) );
BUFX2 BUFX2_1095 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf13_) );
BUFX2 BUFX2_1096 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf12_) );
BUFX2 BUFX2_1097 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf11_) );
BUFX2 BUFX2_1098 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf10_) );
BUFX2 BUFX2_1099 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf9_) );
BUFX2 BUFX2_1100 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf8_) );
BUFX2 BUFX2_1101 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf7_) );
BUFX2 BUFX2_1102 ( .A(decoded_rs1_0__hier0_bF_buf4), .Y(decoded_rs1_0_bF_buf6_) );
BUFX2 BUFX2_1103 ( .A(decoded_rs1_0__hier0_bF_buf3), .Y(decoded_rs1_0_bF_buf5_) );
BUFX2 BUFX2_1104 ( .A(decoded_rs1_0__hier0_bF_buf2), .Y(decoded_rs1_0_bF_buf4_) );
BUFX2 BUFX2_1105 ( .A(decoded_rs1_0__hier0_bF_buf1), .Y(decoded_rs1_0_bF_buf3_) );
BUFX2 BUFX2_1106 ( .A(decoded_rs1_0__hier0_bF_buf0), .Y(decoded_rs1_0_bF_buf2_) );
BUFX2 BUFX2_1107 ( .A(decoded_rs1_0__hier0_bF_buf6), .Y(decoded_rs1_0_bF_buf1_) );
BUFX2 BUFX2_1108 ( .A(decoded_rs1_0__hier0_bF_buf5), .Y(decoded_rs1_0_bF_buf0_) );
BUFX2 BUFX2_1109 ( .A(_4538_), .Y(_4538__bF_buf4) );
BUFX2 BUFX2_1110 ( .A(_4538_), .Y(_4538__bF_buf3) );
BUFX2 BUFX2_1111 ( .A(_4538_), .Y(_4538__bF_buf2) );
BUFX2 BUFX2_1112 ( .A(_4538_), .Y(_4538__bF_buf1) );
BUFX2 BUFX2_1113 ( .A(_4538_), .Y(_4538__bF_buf0) );
BUFX2 BUFX2_1114 ( .A(_3007_), .Y(_3007__bF_buf4) );
BUFX2 BUFX2_1115 ( .A(_3007_), .Y(_3007__bF_buf3) );
BUFX2 BUFX2_1116 ( .A(_3007_), .Y(_3007__bF_buf2) );
BUFX2 BUFX2_1117 ( .A(_3007_), .Y(_3007__bF_buf1) );
BUFX2 BUFX2_1118 ( .A(_3007_), .Y(_3007__bF_buf0) );
BUFX2 BUFX2_1119 ( .A(cpu_state_3_), .Y(cpu_state_3_bF_buf4_) );
BUFX2 BUFX2_1120 ( .A(cpu_state_3_), .Y(cpu_state_3_bF_buf3_) );
BUFX2 BUFX2_1121 ( .A(cpu_state_3_), .Y(cpu_state_3_bF_buf2_) );
BUFX2 BUFX2_1122 ( .A(cpu_state_3_), .Y(cpu_state_3_bF_buf1_) );
BUFX2 BUFX2_1123 ( .A(cpu_state_3_), .Y(cpu_state_3_bF_buf0_) );
BUFX2 BUFX2_1124 ( .A(_10728__1_), .Y(_10728__1_bF_buf3_) );
BUFX2 BUFX2_1125 ( .A(_10728__1_), .Y(_10728__1_bF_buf2_) );
BUFX2 BUFX2_1126 ( .A(_10728__1_), .Y(_10728__1_bF_buf1_) );
BUFX2 BUFX2_1127 ( .A(_10728__1_), .Y(_10728__1_bF_buf0_) );
BUFX2 BUFX2_1128 ( .A(_4632_), .Y(_4632__bF_buf8) );
BUFX2 BUFX2_1129 ( .A(_4632_), .Y(_4632__bF_buf7) );
BUFX2 BUFX2_1130 ( .A(_4632_), .Y(_4632__bF_buf6) );
BUFX2 BUFX2_1131 ( .A(_4632_), .Y(_4632__bF_buf5) );
BUFX2 BUFX2_1132 ( .A(_4632_), .Y(_4632__bF_buf4) );
BUFX2 BUFX2_1133 ( .A(_4632_), .Y(_4632__bF_buf3) );
BUFX2 BUFX2_1134 ( .A(_4632_), .Y(_4632__bF_buf2) );
BUFX2 BUFX2_1135 ( .A(_4632_), .Y(_4632__bF_buf1) );
BUFX2 BUFX2_1136 ( .A(_4632_), .Y(_4632__bF_buf0) );
BUFX2 BUFX2_1137 ( .A(_1566_), .Y(_1566__bF_buf3) );
BUFX2 BUFX2_1138 ( .A(_1566_), .Y(_1566__bF_buf2) );
BUFX2 BUFX2_1139 ( .A(_1566_), .Y(_1566__bF_buf1) );
BUFX2 BUFX2_1140 ( .A(_1566_), .Y(_1566__bF_buf0) );
BUFX2 BUFX2_1141 ( .A(_4917_), .Y(_4917__bF_buf10) );
BUFX2 BUFX2_1142 ( .A(_4917_), .Y(_4917__bF_buf9) );
BUFX2 BUFX2_1143 ( .A(_4917_), .Y(_4917__bF_buf8) );
BUFX2 BUFX2_1144 ( .A(_4917_), .Y(_4917__bF_buf7) );
BUFX2 BUFX2_1145 ( .A(_4917_), .Y(_4917__bF_buf6) );
BUFX2 BUFX2_1146 ( .A(_4917_), .Y(_4917__bF_buf5) );
BUFX2 BUFX2_1147 ( .A(_4917_), .Y(_4917__bF_buf4) );
BUFX2 BUFX2_1148 ( .A(_4917_), .Y(_4917__bF_buf3) );
BUFX2 BUFX2_1149 ( .A(_4917_), .Y(_4917__bF_buf2) );
BUFX2 BUFX2_1150 ( .A(_4917_), .Y(_4917__bF_buf1) );
BUFX2 BUFX2_1151 ( .A(_4917_), .Y(_4917__bF_buf0) );
BUFX2 BUFX2_1152 ( .A(_4955_), .Y(_4955__bF_buf4) );
BUFX2 BUFX2_1153 ( .A(_4955_), .Y(_4955__bF_buf3) );
BUFX2 BUFX2_1154 ( .A(_4955_), .Y(_4955__bF_buf2) );
BUFX2 BUFX2_1155 ( .A(_4955_), .Y(_4955__bF_buf1) );
BUFX2 BUFX2_1156 ( .A(_4955_), .Y(_4955__bF_buf0) );
BUFX2 BUFX2_1157 ( .A(_5358_), .Y(_5358__bF_buf12) );
BUFX2 BUFX2_1158 ( .A(_5358_), .Y(_5358__bF_buf11) );
BUFX2 BUFX2_1159 ( .A(_5358_), .Y(_5358__bF_buf10) );
BUFX2 BUFX2_1160 ( .A(_5358_), .Y(_5358__bF_buf9) );
BUFX2 BUFX2_1161 ( .A(_5358_), .Y(_5358__bF_buf8) );
BUFX2 BUFX2_1162 ( .A(_5358_), .Y(_5358__bF_buf7) );
BUFX2 BUFX2_1163 ( .A(_5358_), .Y(_5358__bF_buf6) );
BUFX2 BUFX2_1164 ( .A(_5358_), .Y(_5358__bF_buf5) );
BUFX2 BUFX2_1165 ( .A(_5358_), .Y(_5358__bF_buf4) );
BUFX2 BUFX2_1166 ( .A(_5358_), .Y(_5358__bF_buf3) );
BUFX2 BUFX2_1167 ( .A(_5358_), .Y(_5358__bF_buf2) );
BUFX2 BUFX2_1168 ( .A(_5358_), .Y(_5358__bF_buf1) );
BUFX2 BUFX2_1169 ( .A(_5358_), .Y(_5358__bF_buf0) );
BUFX2 BUFX2_1170 ( .A(_3844_), .Y(_3844__bF_buf8) );
BUFX2 BUFX2_1171 ( .A(_3844_), .Y(_3844__bF_buf7) );
BUFX2 BUFX2_1172 ( .A(_3844_), .Y(_3844__bF_buf6) );
BUFX2 BUFX2_1173 ( .A(_3844_), .Y(_3844__bF_buf5) );
BUFX2 BUFX2_1174 ( .A(_3844_), .Y(_3844__bF_buf4) );
BUFX2 BUFX2_1175 ( .A(_3844_), .Y(_3844__bF_buf3) );
BUFX2 BUFX2_1176 ( .A(_3844_), .Y(_3844__bF_buf2) );
BUFX2 BUFX2_1177 ( .A(_3844_), .Y(_3844__bF_buf1) );
BUFX2 BUFX2_1178 ( .A(_3844_), .Y(_3844__bF_buf0) );
BUFX2 BUFX2_1179 ( .A(_2313_), .Y(_2313__bF_buf3) );
BUFX2 BUFX2_1180 ( .A(_2313_), .Y(_2313__bF_buf2) );
BUFX2 BUFX2_1181 ( .A(_2313_), .Y(_2313__bF_buf1) );
BUFX2 BUFX2_1182 ( .A(_2313_), .Y(_2313__bF_buf0) );
BUFX2 BUFX2_1183 ( .A(_10103_), .Y(_10103__bF_buf6) );
BUFX2 BUFX2_1184 ( .A(_10103_), .Y(_10103__bF_buf5) );
BUFX2 BUFX2_1185 ( .A(_10103_), .Y(_10103__bF_buf4) );
BUFX2 BUFX2_1186 ( .A(_10103_), .Y(_10103__bF_buf3) );
BUFX2 BUFX2_1187 ( .A(_10103_), .Y(_10103__bF_buf2) );
BUFX2 BUFX2_1188 ( .A(_10103_), .Y(_10103__bF_buf1) );
BUFX2 BUFX2_1189 ( .A(_10103_), .Y(_10103__bF_buf0) );
BUFX2 BUFX2_1190 ( .A(_4664_), .Y(_4664__bF_buf4) );
BUFX2 BUFX2_1191 ( .A(_4664_), .Y(_4664__bF_buf3) );
BUFX2 BUFX2_1192 ( .A(_4664_), .Y(_4664__bF_buf2) );
BUFX2 BUFX2_1193 ( .A(_4664_), .Y(_4664__bF_buf1) );
BUFX2 BUFX2_1194 ( .A(_4664_), .Y(_4664__bF_buf0) );
BUFX2 BUFX2_1195 ( .A(_2310_), .Y(_2310__bF_buf7) );
BUFX2 BUFX2_1196 ( .A(_2310_), .Y(_2310__bF_buf6) );
BUFX2 BUFX2_1197 ( .A(_2310_), .Y(_2310__bF_buf5) );
BUFX2 BUFX2_1198 ( .A(_2310_), .Y(_2310__bF_buf4) );
BUFX2 BUFX2_1199 ( .A(_2310_), .Y(_2310__bF_buf3) );
BUFX2 BUFX2_1200 ( .A(_2310_), .Y(_2310__bF_buf2) );
BUFX2 BUFX2_1201 ( .A(_2310_), .Y(_2310__bF_buf1) );
BUFX2 BUFX2_1202 ( .A(_2310_), .Y(_2310__bF_buf0) );
BUFX2 BUFX2_1203 ( .A(_4893_), .Y(_4893__bF_buf4) );
BUFX2 BUFX2_1204 ( .A(_4893_), .Y(_4893__bF_buf3) );
BUFX2 BUFX2_1205 ( .A(_4893_), .Y(_4893__bF_buf2) );
BUFX2 BUFX2_1206 ( .A(_4893_), .Y(_4893__bF_buf1) );
BUFX2 BUFX2_1207 ( .A(_4893_), .Y(_4893__bF_buf0) );
BUFX2 BUFX2_1208 ( .A(_2345_), .Y(_2345__bF_buf4) );
BUFX2 BUFX2_1209 ( .A(_2345_), .Y(_2345__bF_buf3) );
BUFX2 BUFX2_1210 ( .A(_2345_), .Y(_2345__bF_buf2) );
BUFX2 BUFX2_1211 ( .A(_2345_), .Y(_2345__bF_buf1) );
BUFX2 BUFX2_1212 ( .A(_2345_), .Y(_2345__bF_buf0) );
BUFX2 BUFX2_1213 ( .A(_5314_), .Y(_5314__bF_buf7) );
BUFX2 BUFX2_1214 ( .A(_5314_), .Y(_5314__bF_buf6) );
BUFX2 BUFX2_1215 ( .A(_5314_), .Y(_5314__bF_buf5) );
BUFX2 BUFX2_1216 ( .A(_5314_), .Y(_5314__bF_buf4) );
BUFX2 BUFX2_1217 ( .A(_5314_), .Y(_5314__bF_buf3) );
BUFX2 BUFX2_1218 ( .A(_5314_), .Y(_5314__bF_buf2) );
BUFX2 BUFX2_1219 ( .A(_5314_), .Y(_5314__bF_buf1) );
BUFX2 BUFX2_1220 ( .A(_5314_), .Y(_5314__bF_buf0) );
BUFX2 BUFX2_1221 ( .A(_4755_), .Y(_4755__bF_buf4) );
BUFX2 BUFX2_1222 ( .A(_4755_), .Y(_4755__bF_buf3) );
BUFX2 BUFX2_1223 ( .A(_4755_), .Y(_4755__bF_buf2) );
BUFX2 BUFX2_1224 ( .A(_4755_), .Y(_4755__bF_buf1) );
BUFX2 BUFX2_1225 ( .A(_4755_), .Y(_4755__bF_buf0) );
BUFX2 BUFX2_1226 ( .A(_5349_), .Y(_5349__bF_buf11) );
BUFX2 BUFX2_1227 ( .A(_5349_), .Y(_5349__bF_buf10) );
BUFX2 BUFX2_1228 ( .A(_5349_), .Y(_5349__bF_buf9) );
BUFX2 BUFX2_1229 ( .A(_5349_), .Y(_5349__bF_buf8) );
BUFX2 BUFX2_1230 ( .A(_5349_), .Y(_5349__bF_buf7) );
BUFX2 BUFX2_1231 ( .A(_5349_), .Y(_5349__bF_buf6) );
BUFX2 BUFX2_1232 ( .A(_5349_), .Y(_5349__bF_buf5) );
BUFX2 BUFX2_1233 ( .A(_5349_), .Y(_5349__bF_buf4) );
BUFX2 BUFX2_1234 ( .A(_5349_), .Y(_5349__bF_buf3) );
BUFX2 BUFX2_1235 ( .A(_5349_), .Y(_5349__bF_buf2) );
BUFX2 BUFX2_1236 ( .A(_5349_), .Y(_5349__bF_buf1) );
BUFX2 BUFX2_1237 ( .A(_5349_), .Y(_5349__bF_buf0) );
BUFX2 BUFX2_1238 ( .A(_4793_), .Y(_4793__bF_buf4) );
BUFX2 BUFX2_1239 ( .A(_4793_), .Y(_4793__bF_buf3) );
BUFX2 BUFX2_1240 ( .A(_4793_), .Y(_4793__bF_buf2) );
BUFX2 BUFX2_1241 ( .A(_4793_), .Y(_4793__bF_buf1) );
BUFX2 BUFX2_1242 ( .A(_4793_), .Y(_4793__bF_buf0) );
BUFX2 BUFX2_1243 ( .A(_4047_), .Y(_4047__bF_buf7) );
BUFX2 BUFX2_1244 ( .A(_4047_), .Y(_4047__bF_buf6) );
BUFX2 BUFX2_1245 ( .A(_4047_), .Y(_4047__bF_buf5) );
BUFX2 BUFX2_1246 ( .A(_4047_), .Y(_4047__bF_buf4) );
BUFX2 BUFX2_1247 ( .A(_4047_), .Y(_4047__bF_buf3) );
BUFX2 BUFX2_1248 ( .A(_4047_), .Y(_4047__bF_buf2) );
BUFX2 BUFX2_1249 ( .A(_4047_), .Y(_4047__bF_buf1) );
BUFX2 BUFX2_1250 ( .A(_4047_), .Y(_4047__bF_buf0) );
BUFX2 BUFX2_1251 ( .A(_4696_), .Y(_4696__bF_buf4) );
BUFX2 BUFX2_1252 ( .A(_4696_), .Y(_4696__bF_buf3) );
BUFX2 BUFX2_1253 ( .A(_4696_), .Y(_4696__bF_buf2) );
BUFX2 BUFX2_1254 ( .A(_4696_), .Y(_4696__bF_buf1) );
BUFX2 BUFX2_1255 ( .A(_4696_), .Y(_4696__bF_buf0) );
BUFX2 BUFX2_1256 ( .A(_3776_), .Y(_3776__bF_buf7) );
BUFX2 BUFX2_1257 ( .A(_3776_), .Y(_3776__bF_buf6) );
BUFX2 BUFX2_1258 ( .A(_3776_), .Y(_3776__bF_buf5) );
BUFX2 BUFX2_1259 ( .A(_3776_), .Y(_3776__bF_buf4) );
BUFX2 BUFX2_1260 ( .A(_3776_), .Y(_3776__bF_buf3) );
BUFX2 BUFX2_1261 ( .A(_3776_), .Y(_3776__bF_buf2) );
BUFX2 BUFX2_1262 ( .A(_3776_), .Y(_3776__bF_buf1) );
BUFX2 BUFX2_1263 ( .A(_3776_), .Y(_3776__bF_buf0) );
BUFX2 BUFX2_1264 ( .A(_2207_), .Y(_2207__bF_buf4) );
BUFX2 BUFX2_1265 ( .A(_2207_), .Y(_2207__bF_buf3) );
BUFX2 BUFX2_1266 ( .A(_2207_), .Y(_2207__bF_buf2) );
BUFX2 BUFX2_1267 ( .A(_2207_), .Y(_2207__bF_buf1) );
BUFX2 BUFX2_1268 ( .A(_2207_), .Y(_2207__bF_buf0) );
BUFX2 BUFX2_1269 ( .A(_4714_), .Y(_4714__bF_buf3) );
BUFX2 BUFX2_1270 ( .A(_4714_), .Y(_4714__bF_buf2) );
BUFX2 BUFX2_1271 ( .A(_4714_), .Y(_4714__bF_buf1) );
BUFX2 BUFX2_1272 ( .A(_4714_), .Y(_4714__bF_buf0) );
BUFX2 BUFX2_1273 ( .A(_5290_), .Y(_5290__bF_buf3) );
BUFX2 BUFX2_1274 ( .A(_5290_), .Y(_5290__bF_buf2) );
BUFX2 BUFX2_1275 ( .A(_5290_), .Y(_5290__bF_buf1) );
BUFX2 BUFX2_1276 ( .A(_5290_), .Y(_5290__bF_buf0) );
BUFX2 BUFX2_1277 ( .A(_4426_), .Y(_4426__bF_buf11) );
BUFX2 BUFX2_1278 ( .A(_4426_), .Y(_4426__bF_buf10) );
BUFX2 BUFX2_1279 ( .A(_4426_), .Y(_4426__bF_buf9) );
BUFX2 BUFX2_1280 ( .A(_4426_), .Y(_4426__bF_buf8) );
BUFX2 BUFX2_1281 ( .A(_4426_), .Y(_4426__bF_buf7) );
BUFX2 BUFX2_1282 ( .A(_4426_), .Y(_4426__bF_buf6) );
BUFX2 BUFX2_1283 ( .A(_4426_), .Y(_4426__bF_buf5) );
BUFX2 BUFX2_1284 ( .A(_4426_), .Y(_4426__bF_buf4) );
BUFX2 BUFX2_1285 ( .A(_4426_), .Y(_4426__bF_buf3) );
BUFX2 BUFX2_1286 ( .A(_4426_), .Y(_4426__bF_buf2) );
BUFX2 BUFX2_1287 ( .A(_4426_), .Y(_4426__bF_buf1) );
BUFX2 BUFX2_1288 ( .A(_4426_), .Y(_4426__bF_buf0) );
BUFX2 BUFX2_1289 ( .A(_4884_), .Y(_4884__bF_buf4) );
BUFX2 BUFX2_1290 ( .A(_4884_), .Y(_4884__bF_buf3) );
BUFX2 BUFX2_1291 ( .A(_4884_), .Y(_4884__bF_buf2) );
BUFX2 BUFX2_1292 ( .A(_4884_), .Y(_4884__bF_buf1) );
BUFX2 BUFX2_1293 ( .A(_4884_), .Y(_4884__bF_buf0) );
BUFX2 BUFX2_1294 ( .A(_7624_), .Y(_7624__bF_buf4) );
BUFX2 BUFX2_1295 ( .A(_7624_), .Y(_7624__bF_buf3) );
BUFX2 BUFX2_1296 ( .A(_7624_), .Y(_7624__bF_buf2) );
BUFX2 BUFX2_1297 ( .A(_7624_), .Y(_7624__bF_buf1) );
BUFX2 BUFX2_1298 ( .A(_7624_), .Y(_7624__bF_buf0) );
BUFX2 BUFX2_1299 ( .A(_4499_), .Y(_4499__bF_buf5) );
BUFX2 BUFX2_1300 ( .A(_4499_), .Y(_4499__bF_buf4) );
BUFX2 BUFX2_1301 ( .A(_4499_), .Y(_4499__bF_buf3) );
BUFX2 BUFX2_1302 ( .A(_4499_), .Y(_4499__bF_buf2) );
BUFX2 BUFX2_1303 ( .A(_4499_), .Y(_4499__bF_buf1) );
BUFX2 BUFX2_1304 ( .A(_4499_), .Y(_4499__bF_buf0) );
BUFX2 BUFX2_1305 ( .A(_4940_), .Y(_4940__bF_buf4) );
BUFX2 BUFX2_1306 ( .A(_4940_), .Y(_4940__bF_buf3) );
BUFX2 BUFX2_1307 ( .A(_4940_), .Y(_4940__bF_buf2) );
BUFX2 BUFX2_1308 ( .A(_4940_), .Y(_4940__bF_buf1) );
BUFX2 BUFX2_1309 ( .A(_4940_), .Y(_4940__bF_buf0) );
BUFX2 BUFX2_1310 ( .A(_7697_), .Y(_7697__bF_buf3) );
BUFX2 BUFX2_1311 ( .A(_7697_), .Y(_7697__bF_buf2) );
BUFX2 BUFX2_1312 ( .A(_7697_), .Y(_7697__bF_buf1) );
BUFX2 BUFX2_1313 ( .A(_7697_), .Y(_7697__bF_buf0) );
BUFX2 BUFX2_1314 ( .A(_2104_), .Y(_2104__bF_buf7) );
BUFX2 BUFX2_1315 ( .A(_2104_), .Y(_2104__bF_buf6) );
BUFX2 BUFX2_1316 ( .A(_2104_), .Y(_2104__bF_buf5) );
BUFX2 BUFX2_1317 ( .A(_2104_), .Y(_2104__bF_buf4) );
BUFX2 BUFX2_1318 ( .A(_2104_), .Y(_2104__bF_buf3) );
BUFX2 BUFX2_1319 ( .A(_2104_), .Y(_2104__bF_buf2) );
BUFX2 BUFX2_1320 ( .A(_2104_), .Y(_2104__bF_buf1) );
BUFX2 BUFX2_1321 ( .A(_2104_), .Y(_2104__bF_buf0) );
BUFX2 BUFX2_1322 ( .A(_10123_), .Y(_10123__bF_buf4) );
BUFX2 BUFX2_1323 ( .A(_10123_), .Y(_10123__bF_buf3) );
BUFX2 BUFX2_1324 ( .A(_10123_), .Y(_10123__bF_buf2) );
BUFX2 BUFX2_1325 ( .A(_10123_), .Y(_10123__bF_buf1) );
BUFX2 BUFX2_1326 ( .A(_10123_), .Y(_10123__bF_buf0) );
BUFX2 BUFX2_1327 ( .A(_2274_), .Y(_2274__bF_buf4) );
BUFX2 BUFX2_1328 ( .A(_2274_), .Y(_2274__bF_buf3) );
BUFX2 BUFX2_1329 ( .A(_2274_), .Y(_2274__bF_buf2) );
BUFX2 BUFX2_1330 ( .A(_2274_), .Y(_2274__bF_buf1) );
BUFX2 BUFX2_1331 ( .A(_2274_), .Y(_2274__bF_buf0) );
BUFX2 BUFX2_1332 ( .A(_5281_), .Y(_5281__bF_buf10) );
BUFX2 BUFX2_1333 ( .A(_5281_), .Y(_5281__bF_buf9) );
BUFX2 BUFX2_1334 ( .A(_5281_), .Y(_5281__bF_buf8) );
BUFX2 BUFX2_1335 ( .A(_5281_), .Y(_5281__bF_buf7) );
BUFX2 BUFX2_1336 ( .A(_5281_), .Y(_5281__bF_buf6) );
BUFX2 BUFX2_1337 ( .A(_5281_), .Y(_5281__bF_buf5) );
BUFX2 BUFX2_1338 ( .A(_5281_), .Y(_5281__bF_buf4) );
BUFX2 BUFX2_1339 ( .A(_5281_), .Y(_5281__bF_buf3) );
BUFX2 BUFX2_1340 ( .A(_5281_), .Y(_5281__bF_buf2) );
BUFX2 BUFX2_1341 ( .A(_5281_), .Y(_5281__bF_buf1) );
BUFX2 BUFX2_1342 ( .A(_5281_), .Y(_5281__bF_buf0) );
INVX1 INVX1_1 ( .A(mem_wordsize_0_bF_buf3_), .Y(_4425_) );
INVX1 INVX1_2 ( .A(resetn_bF_buf11), .Y(_4426_) );
INVX1 INVX1_3 ( .A(mem_do_rdata), .Y(_4427_) );
NOR2X1 NOR2X1_1 ( .A(_4426__bF_buf11), .B(_4427_), .Y(_4428_) );
INVX1 INVX1_4 ( .A(_4428_), .Y(_4429_) );
INVX1 INVX1_5 ( .A(mem_do_prefetch_bF_buf5), .Y(_4430_) );
INVX1 INVX1_6 ( .A(cpu_state_1_bF_buf5_), .Y(_4431_) );
INVX1 INVX1_7 ( .A(mem_state_1_), .Y(_4432_) );
INVX1 INVX1_8 ( .A(mem_state_0_), .Y(_4433_) );
NOR2X1 NOR2X1_2 ( .A(_4432_), .B(_4433_), .Y(_4434_) );
INVX1 INVX1_9 ( .A(mem_do_wdata), .Y(_4435_) );
NOR2X1 NOR2X1_3 ( .A(mem_do_rinst_bF_buf4), .B(mem_do_rdata), .Y(_4436_) );
NAND2X1 NAND2X1_1 ( .A(_4435_), .B(_4436_), .Y(_4437_) );
NOR2X1 NOR2X1_4 ( .A(mem_state_1_), .B(mem_state_0_), .Y(_4438_) );
NAND2X1 NAND2X1_2 ( .A(mem_ready), .B(_10731_), .Y(_4439_) );
NOR2X1 NOR2X1_5 ( .A(_4439__bF_buf6), .B(_4438_), .Y(_4440_) );
AOI22X1 AOI22X1_1 ( .A(mem_do_rinst_bF_buf3), .B(_4434_), .C(_4440_), .D(_4437_), .Y(_4441_) );
NOR2X1 NOR2X1_6 ( .A(_4426__bF_buf10), .B(_4441_), .Y(_4442_) );
OAI21X1 OAI21X1_1 ( .A(_4442_), .B(_4430_), .C(_4431__bF_buf7), .Y(_4443_) );
INVX1 INVX1_10 ( .A(_4443_), .Y(_4444_) );
NOR2X1 NOR2X1_7 ( .A(cpu_state_4_), .B(cpu_state_2_bF_buf5_), .Y(_4445_) );
INVX1 INVX1_11 ( .A(_4445_), .Y(_4446_) );
NOR2X1 NOR2X1_8 ( .A(cpu_state_3_bF_buf4_), .B(_4446_), .Y(_4447_) );
INVX1 INVX1_12 ( .A(_4447__bF_buf3), .Y(_4448_) );
NOR2X1 NOR2X1_9 ( .A(cpu_state_5_bF_buf3_), .B(cpu_state_0_), .Y(_4449_) );
INVX1 INVX1_13 ( .A(_4449_), .Y(_4450_) );
NOR2X1 NOR2X1_10 ( .A(_4450_), .B(_4448_), .Y(_4451_) );
NAND2X1 NAND2X1_3 ( .A(_4451_), .B(_4444_), .Y(_4452_) );
OAI21X1 OAI21X1_2 ( .A(_4441_), .B(_4426__bF_buf9), .C(mem_do_prefetch_bF_buf4), .Y(_4453_) );
INVX1 INVX1_14 ( .A(_4453_), .Y(_4454_) );
NAND2X1 NAND2X1_4 ( .A(resetn_bF_buf10), .B(_4441_), .Y(_4455_) );
INVX1 INVX1_15 ( .A(_4455_), .Y(_4456_) );
NAND2X1 NAND2X1_5 ( .A(mem_do_prefetch_bF_buf3), .B(_4456_), .Y(_4457_) );
NOR2X1 NOR2X1_11 ( .A(_4426__bF_buf8), .B(_4435_), .Y(_4458_) );
INVX1 INVX1_16 ( .A(_4458_), .Y(_4459_) );
OAI21X1 OAI21X1_3 ( .A(_4454_), .B(_4459_), .C(_4457_), .Y(_4460_) );
NOR2X1 NOR2X1_12 ( .A(cpu_state_5_bF_buf2_), .B(cpu_state_1_bF_buf4_), .Y(_4461_) );
NOR2X1 NOR2X1_13 ( .A(cpu_state_0_), .B(_4426__bF_buf7), .Y(_4462_) );
NAND2X1 NAND2X1_6 ( .A(_4462_), .B(_4447__bF_buf2), .Y(_4463_) );
AOI21X1 AOI21X1_1 ( .A(_4461_), .B(_4454_), .C(_4463_), .Y(_4464_) );
INVX1 INVX1_17 ( .A(_4464_), .Y(_4465_) );
AOI21X1 AOI21X1_2 ( .A(cpu_state_5_bF_buf1_), .B(_4460_), .C(_4465_), .Y(_4466_) );
OAI21X1 OAI21X1_4 ( .A(_4429_), .B(_4452_), .C(_4466_), .Y(_4467_) );
INVX1 INVX1_18 ( .A(_4467_), .Y(_4468_) );
NOR2X1 NOR2X1_14 ( .A(instr_sh), .B(instr_sb), .Y(_4469_) );
NAND2X1 NAND2X1_7 ( .A(cpu_state_5_bF_buf0_), .B(_4435_), .Y(_4470_) );
OAI21X1 OAI21X1_5 ( .A(_4442_), .B(_4430_), .C(resetn_bF_buf9), .Y(_4471_) );
NOR2X1 NOR2X1_15 ( .A(_4470_), .B(_4471_), .Y(_4472_) );
NAND2X1 NAND2X1_8 ( .A(_4469_), .B(_4472_), .Y(_4473_) );
NOR2X1 NOR2X1_16 ( .A(_4426__bF_buf6), .B(_4431__bF_buf6), .Y(_4474_) );
INVX1 INVX1_19 ( .A(_4474_), .Y(_4475_) );
NOR2X1 NOR2X1_17 ( .A(mem_do_rdata), .B(_4426__bF_buf5), .Y(_4476_) );
NOR2X1 NOR2X1_18 ( .A(instr_lh), .B(instr_lb), .Y(_4477_) );
NOR2X1 NOR2X1_19 ( .A(instr_lhu), .B(instr_lbu), .Y(_4478_) );
AND2X2 AND2X2_1 ( .A(_4477_), .B(_4478_), .Y(_4479_) );
AND2X2 AND2X2_2 ( .A(_4451_), .B(_4479_), .Y(_4480_) );
NAND3X1 NAND3X1_1 ( .A(_4476_), .B(_4480_), .C(_4444_), .Y(_4481_) );
NAND3X1 NAND3X1_2 ( .A(_4475_), .B(_4481_), .C(_4473_), .Y(_4482_) );
INVX1 INVX1_20 ( .A(_4482_), .Y(_4483_) );
OAI21X1 OAI21X1_6 ( .A(_4468_), .B(_4425_), .C(_4483_), .Y(_378_) );
OAI21X1 OAI21X1_7 ( .A(instr_lh), .B(instr_lhu), .C(_4476_), .Y(_4484_) );
AOI22X1 AOI22X1_2 ( .A(instr_sh), .B(_4472_), .C(_4467_), .D(mem_wordsize_2_), .Y(_4485_) );
OAI21X1 OAI21X1_8 ( .A(_4452_), .B(_4484_), .C(_4485_), .Y(_87_) );
OAI21X1 OAI21X1_9 ( .A(reg_pc_0_), .B(reg_pc_1_), .C(mem_do_rinst_bF_buf2), .Y(_4486_) );
NOR2X1 NOR2X1_20 ( .A(_4426__bF_buf4), .B(_4486_), .Y(_4487_) );
INVX1 INVX1_21 ( .A(_4487_), .Y(_4488_) );
OAI21X1 OAI21X1_10 ( .A(mem_do_wdata), .B(mem_do_rdata), .C(resetn_bF_buf8), .Y(_4489_) );
INVX1 INVX1_22 ( .A(_10734__1_), .Y(_4490_) );
INVX1 INVX1_23 ( .A(_10734__0_), .Y(_4491_) );
OAI21X1 OAI21X1_11 ( .A(_4425_), .B(_4490_), .C(_4491_), .Y(_4492_) );
OAI21X1 OAI21X1_12 ( .A(mem_wordsize_0_bF_buf2_), .B(mem_wordsize_2_), .C(_4492_), .Y(_4493_) );
OAI21X1 OAI21X1_13 ( .A(_4493_), .B(_4489_), .C(_4488_), .Y(_4494_) );
INVX1 INVX1_24 ( .A(_4489_), .Y(_4495_) );
OAI21X1 OAI21X1_14 ( .A(_4428_), .B(_4458_), .C(_4493_), .Y(_4496_) );
OAI21X1 OAI21X1_15 ( .A(_4426__bF_buf3), .B(_4495_), .C(_4496_), .Y(_4497_) );
AOI21X1 AOI21X1_3 ( .A(cpu_state_0_), .B(_4497_), .C(_4494_), .Y(_4498_) );
INVX1 INVX1_25 ( .A(instr_jal_bF_buf6), .Y(_4499_) );
NOR2X1 NOR2X1_21 ( .A(instr_lui), .B(instr_auipc), .Y(_4500_) );
NAND2X1 NAND2X1_9 ( .A(_4499__bF_buf5), .B(_4500_), .Y(_57_) );
NOR2X1 NOR2X1_22 ( .A(instr_slti), .B(instr_slt), .Y(_4501_) );
NOR2X1 NOR2X1_23 ( .A(instr_sltiu), .B(instr_sltu), .Y(_4502_) );
NAND2X1 NAND2X1_10 ( .A(_4501_), .B(_4502_), .Y(_4503_) );
NOR2X1 NOR2X1_24 ( .A(_57_), .B(_4503_), .Y(_4504_) );
NOR2X1 NOR2X1_25 ( .A(instr_bgeu), .B(instr_beq), .Y(_4505_) );
NOR2X1 NOR2X1_26 ( .A(instr_bge), .B(instr_bne), .Y(_4506_) );
NAND2X1 NAND2X1_11 ( .A(_4505_), .B(_4506_), .Y(_4507_) );
NOR2X1 NOR2X1_27 ( .A(instr_add), .B(instr_sub_bF_buf4), .Y(_4508_) );
NOR2X1 NOR2X1_28 ( .A(instr_jalr), .B(instr_addi), .Y(_4509_) );
NAND2X1 NAND2X1_12 ( .A(_4508_), .B(_4509_), .Y(_4510_) );
NOR2X1 NOR2X1_29 ( .A(_4510_), .B(_4507_), .Y(_4511_) );
NAND2X1 NAND2X1_13 ( .A(_4504_), .B(_4511_), .Y(_4512_) );
NOR2X1 NOR2X1_30 ( .A(instr_or), .B(instr_and), .Y(_4513_) );
NOR2X1 NOR2X1_31 ( .A(instr_srl), .B(instr_sra), .Y(_4514_) );
NAND2X1 NAND2X1_14 ( .A(_4513_), .B(_4514_), .Y(_4515_) );
INVX1 INVX1_26 ( .A(instr_srli), .Y(_4516_) );
INVX1 INVX1_27 ( .A(instr_srai), .Y(_4517_) );
NOR2X1 NOR2X1_32 ( .A(instr_sll), .B(instr_xor), .Y(_4518_) );
NAND3X1 NAND3X1_3 ( .A(_4516_), .B(_4517_), .C(_4518_), .Y(_4519_) );
NOR2X1 NOR2X1_33 ( .A(_4515_), .B(_4519_), .Y(_4520_) );
INVX1 INVX1_28 ( .A(instr_lw), .Y(_4521_) );
INVX1 INVX1_29 ( .A(instr_blt), .Y(_4522_) );
NOR2X1 NOR2X1_34 ( .A(instr_xori), .B(instr_ori), .Y(_4523_) );
NAND3X1 NAND3X1_4 ( .A(_4521_), .B(_4522_), .C(_4523_), .Y(_4524_) );
NOR2X1 NOR2X1_35 ( .A(instr_andi), .B(instr_slli), .Y(_4525_) );
NOR2X1 NOR2X1_36 ( .A(instr_sw), .B(instr_bltu), .Y(_4526_) );
NAND2X1 NAND2X1_15 ( .A(_4525_), .B(_4526_), .Y(_4527_) );
NOR2X1 NOR2X1_37 ( .A(_4527_), .B(_4524_), .Y(_4528_) );
INVX1 INVX1_30 ( .A(instr_rdinstr_bF_buf4), .Y(_4529_) );
NOR2X1 NOR2X1_38 ( .A(instr_rdcycle_bF_buf4), .B(instr_rdcycleh_bF_buf3), .Y(_4530_) );
NAND2X1 NAND2X1_16 ( .A(_4529_), .B(_4530_), .Y(_4531_) );
NOR2X1 NOR2X1_39 ( .A(instr_rdinstrh), .B(_4531__bF_buf4), .Y(_4532_) );
INVX1 INVX1_31 ( .A(_4532_), .Y(_4533_) );
NAND3X1 NAND3X1_5 ( .A(_4469_), .B(_4477_), .C(_4478_), .Y(_4534_) );
NOR2X1 NOR2X1_40 ( .A(_4534_), .B(_4533_), .Y(_4535_) );
NAND3X1 NAND3X1_6 ( .A(_4520_), .B(_4528_), .C(_4535_), .Y(_4536_) );
OR2X2 OR2X2_1 ( .A(_4536_), .B(_4512_), .Y(_4537_) );
INVX1 INVX1_32 ( .A(cpu_state_2_bF_buf4_), .Y(_4538_) );
NOR2X1 NOR2X1_41 ( .A(_4426__bF_buf2), .B(_4538__bF_buf4), .Y(_4539_) );
INVX1 INVX1_33 ( .A(_4539__bF_buf3), .Y(_4540_) );
OAI21X1 OAI21X1_16 ( .A(_4537_), .B(_4540__bF_buf6), .C(_4498_), .Y(_88_) );
NAND2X1 NAND2X1_17 ( .A(_4522_), .B(_4501_), .Y(_62_) );
NAND2X1 NAND2X1_18 ( .A(_4521_), .B(_4478_), .Y(_56_) );
INVX1 INVX1_34 ( .A(mem_rdata_q_3_), .Y(_4541_) );
INVX1 INVX1_35 ( .A(_4439__bF_buf5), .Y(_4542_) );
NAND2X1 NAND2X1_19 ( .A(mem_rdata[3]), .B(_4542_), .Y(_4543_) );
OAI21X1 OAI21X1_17 ( .A(_4541_), .B(_4542_), .C(_4543_), .Y(mem_rdata_latched_3_) );
INVX1 INVX1_36 ( .A(mem_rdata[4]), .Y(_4544_) );
NAND2X1 NAND2X1_20 ( .A(mem_rdata_q_4_), .B(_4439__bF_buf4), .Y(_4545_) );
OAI21X1 OAI21X1_18 ( .A(_4544_), .B(_4439__bF_buf3), .C(_4545_), .Y(mem_rdata_latched_4_) );
INVX1 INVX1_37 ( .A(mem_rdata_q_5_), .Y(_4546_) );
NAND2X1 NAND2X1_21 ( .A(mem_rdata[5]), .B(_4542_), .Y(_4547_) );
OAI21X1 OAI21X1_19 ( .A(_4546_), .B(_4542_), .C(_4547_), .Y(mem_rdata_latched_5_) );
MUX2X1 MUX2X1_1 ( .A(mem_rdata_q_6_), .B(mem_rdata[6]), .S(_4439__bF_buf2), .Y(_4548_) );
INVX1 INVX1_38 ( .A(_4548_), .Y(mem_rdata_latched_6_) );
INVX1 INVX1_39 ( .A(mem_rdata[2]), .Y(_4549_) );
NAND2X1 NAND2X1_22 ( .A(mem_rdata_q_2_), .B(_4439__bF_buf1), .Y(_4550_) );
OAI21X1 OAI21X1_20 ( .A(_4549_), .B(_4439__bF_buf0), .C(_4550_), .Y(mem_rdata_latched_2_) );
INVX1 INVX1_40 ( .A(_4494_), .Y(_4551_) );
NOR2X1 NOR2X1_42 ( .A(is_lui_auipc_jal), .B(is_jalr_addi_slti_sltiu_xori_ori_andi), .Y(_4552_) );
NOR2X1 NOR2X1_43 ( .A(_4538__bF_buf3), .B(_4552_), .Y(_4553_) );
AND2X2 AND2X2_3 ( .A(_4488_), .B(_4553_), .Y(_4554_) );
INVX1 INVX1_41 ( .A(cpu_state_3_bF_buf3_), .Y(_4555_) );
INVX1 INVX1_42 ( .A(is_beq_bne_blt_bge_bltu_bgeu), .Y(_4556_) );
NOR2X1 NOR2X1_44 ( .A(_4555_), .B(_4556_), .Y(_4557_) );
INVX1 INVX1_43 ( .A(_4557_), .Y(_4558_) );
NOR2X1 NOR2X1_45 ( .A(_4558_), .B(_4455_), .Y(_4559_) );
AOI22X1 AOI22X1_3 ( .A(_4497_), .B(_4554_), .C(_4559_), .D(_4551_), .Y(_4560_) );
OAI21X1 OAI21X1_21 ( .A(_4536_), .B(_4512_), .C(_4532_), .Y(_4561_) );
NOR2X1 NOR2X1_46 ( .A(_4426__bF_buf1), .B(_4561_), .Y(_4562_) );
INVX1 INVX1_44 ( .A(_4562_), .Y(_4563_) );
INVX1 INVX1_45 ( .A(is_slli_srli_srai), .Y(_4564_) );
OAI21X1 OAI21X1_22 ( .A(_4536_), .B(_4512_), .C(is_lb_lh_lw_lbu_lhu), .Y(_4565_) );
AND2X2 AND2X2_4 ( .A(_4565_), .B(_4564_), .Y(_4566_) );
NAND2X1 NAND2X1_23 ( .A(cpu_state_2_bF_buf3_), .B(_4552_), .Y(_4567_) );
NOR2X1 NOR2X1_47 ( .A(is_sb_sh_sw), .B(is_sll_srl_sra), .Y(_4568_) );
INVX1 INVX1_46 ( .A(_4568_), .Y(_4569_) );
NOR2X1 NOR2X1_48 ( .A(_4569_), .B(_4567_), .Y(_4570_) );
NAND3X1 NAND3X1_7 ( .A(_4551_), .B(_4570_), .C(_4566_), .Y(_4571_) );
OAI21X1 OAI21X1_23 ( .A(_4571_), .B(_4563_), .C(_4560_), .Y(_89_) );
INVX1 INVX1_47 ( .A(is_sll_srl_sra), .Y(_4572_) );
NOR2X1 NOR2X1_49 ( .A(_4572_), .B(_4567_), .Y(_4573_) );
NAND3X1 NAND3X1_8 ( .A(_4562_), .B(_4573_), .C(_4566_), .Y(_4574_) );
INVX1 INVX1_48 ( .A(cpu_state_4_), .Y(_4575_) );
INVX1 INVX1_49 ( .A(reg_sh_1_), .Y(_4576_) );
NOR2X1 NOR2X1_50 ( .A(reg_sh_3_), .B(reg_sh_2_), .Y(_4577_) );
INVX1 INVX1_50 ( .A(_4577_), .Y(_4578_) );
NOR2X1 NOR2X1_51 ( .A(reg_sh_4_), .B(_4578_), .Y(_4579_) );
INVX1 INVX1_51 ( .A(_4579__bF_buf4), .Y(_4580_) );
NOR2X1 NOR2X1_52 ( .A(reg_sh_0_), .B(_4580__bF_buf4), .Y(_4581_) );
NAND2X1 NAND2X1_24 ( .A(_4576_), .B(_4581_), .Y(_4582_) );
INVX1 INVX1_52 ( .A(_4582_), .Y(_4583_) );
NOR2X1 NOR2X1_53 ( .A(_4575__bF_buf4), .B(_4583_), .Y(_4584_) );
NOR2X1 NOR2X1_54 ( .A(_4538__bF_buf2), .B(_4564_), .Y(_4585_) );
OAI21X1 OAI21X1_24 ( .A(_4584_), .B(_4585_), .C(resetn_bF_buf7), .Y(_4586_) );
AOI21X1 AOI21X1_4 ( .A(_4586_), .B(_4574_), .C(_4494_), .Y(_90_) );
INVX1 INVX1_53 ( .A(cpu_state_5_bF_buf3_), .Y(_4587_) );
INVX1 INVX1_54 ( .A(_4442_), .Y(_4588_) );
NOR2X1 NOR2X1_55 ( .A(mem_do_prefetch_bF_buf2), .B(_4588_), .Y(_4589_) );
OAI21X1 OAI21X1_25 ( .A(_4589_), .B(_4471_), .C(_4457_), .Y(_4590_) );
NAND2X1 NAND2X1_25 ( .A(_4551_), .B(_4590_), .Y(_4591_) );
INVX1 INVX1_55 ( .A(is_sb_sh_sw), .Y(_4592_) );
NOR2X1 NOR2X1_56 ( .A(_4592_), .B(_4567_), .Y(_4593_) );
NAND3X1 NAND3X1_9 ( .A(_4551_), .B(_4593_), .C(_4566_), .Y(_4594_) );
OAI22X1 OAI22X1_1 ( .A(_4587__bF_buf3), .B(_4591_), .C(_4594_), .D(_4563_), .Y(_91_) );
INVX1 INVX1_56 ( .A(cpu_state_6_), .Y(_4595_) );
NAND2X1 NAND2X1_26 ( .A(_4539__bF_buf2), .B(_4551_), .Y(_4596_) );
OAI22X1 OAI22X1_2 ( .A(_4596_), .B(_4565_), .C(_4591_), .D(_4595_), .Y(_92_) );
NOR2X1 NOR2X1_57 ( .A(_4575__bF_buf3), .B(_4582_), .Y(_4597_) );
OAI21X1 OAI21X1_26 ( .A(cpu_state_5_bF_buf2_), .B(cpu_state_6_), .C(_4430_), .Y(_4598_) );
AOI21X1 AOI21X1_5 ( .A(_4558_), .B(_4598_), .C(_4441_), .Y(_4599_) );
OAI21X1 OAI21X1_27 ( .A(_4597__bF_buf3), .B(_4599_), .C(_4551_), .Y(_4600_) );
NOR2X1 NOR2X1_58 ( .A(_4538__bF_buf1), .B(_4532_), .Y(_4601_) );
NOR2X1 NOR2X1_59 ( .A(_4489_), .B(_4493_), .Y(_4602_) );
NAND2X1 NAND2X1_27 ( .A(resetn_bF_buf6), .B(cpu_state_3_bF_buf2_), .Y(_4603_) );
NOR2X1 NOR2X1_60 ( .A(is_beq_bne_blt_bge_bltu_bgeu), .B(_4603_), .Y(_4604_) );
INVX1 INVX1_57 ( .A(decoder_trigger_bF_buf3), .Y(_4605_) );
NOR2X1 NOR2X1_61 ( .A(instr_jal_bF_buf5), .B(_4605__bF_buf5), .Y(_4606_) );
NOR2X1 NOR2X1_62 ( .A(_4431__bF_buf5), .B(_4606_), .Y(_4607_) );
OAI21X1 OAI21X1_28 ( .A(_4607_), .B(_4604_), .C(_4486_), .Y(_4608_) );
OAI21X1 OAI21X1_29 ( .A(_4608_), .B(_4602_), .C(resetn_bF_buf5), .Y(_4609_) );
AOI21X1 AOI21X1_6 ( .A(_4551_), .B(_4601_), .C(_4609_), .Y(_4610_) );
NAND2X1 NAND2X1_28 ( .A(_4610_), .B(_4600_), .Y(_93_) );
INVX1 INVX1_58 ( .A(_4606_), .Y(_4611_) );
NOR2X1 NOR2X1_63 ( .A(_4611_), .B(_4475_), .Y(_4612_) );
AND2X2 AND2X2_5 ( .A(_4551_), .B(_4612_), .Y(_94_) );
INVX1 INVX1_59 ( .A(mem_rdata[12]), .Y(_4613_) );
NAND2X1 NAND2X1_29 ( .A(mem_rdata_q_12_), .B(_4439__bF_buf6), .Y(_4614_) );
OAI21X1 OAI21X1_30 ( .A(_4613_), .B(_4439__bF_buf5), .C(_4614_), .Y(mem_rdata_latched_12_) );
INVX1 INVX1_60 ( .A(mem_rdata[13]), .Y(_4615_) );
NAND2X1 NAND2X1_30 ( .A(mem_rdata_q_13_), .B(_4439__bF_buf4), .Y(_4616_) );
OAI21X1 OAI21X1_31 ( .A(_4615_), .B(_4439__bF_buf3), .C(_4616_), .Y(mem_rdata_latched_13_) );
INVX1 INVX1_61 ( .A(mem_rdata[14]), .Y(_4617_) );
NAND2X1 NAND2X1_31 ( .A(mem_rdata_q_14_), .B(_4439__bF_buf2), .Y(_4618_) );
OAI21X1 OAI21X1_32 ( .A(_4617_), .B(_4439__bF_buf1), .C(_4618_), .Y(mem_rdata_latched_14_) );
INVX1 INVX1_62 ( .A(_4438_), .Y(_4619_) );
NOR2X1 NOR2X1_64 ( .A(_4619_), .B(_4459_), .Y(_10729_) );
NOR2X1 NOR2X1_65 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf1), .Y(_4620_) );
INVX1 INVX1_63 ( .A(_4620_), .Y(_4621_) );
OAI21X1 OAI21X1_33 ( .A(_4621__bF_buf4), .B(mem_do_rdata), .C(_4438_), .Y(_4622_) );
NOR2X1 NOR2X1_66 ( .A(_4426__bF_buf0), .B(_4622_), .Y(_10727_) );
INVX1 INVX1_64 ( .A(cpuregs_8_[5]), .Y(_4623_) );
NOR2X1 NOR2X1_67 ( .A(latched_rd_1_), .B(latched_rd_0_), .Y(_4624_) );
NOR2X1 NOR2X1_68 ( .A(latched_rd_3_), .B(latched_rd_4_), .Y(_4625_) );
INVX1 INVX1_65 ( .A(_4625_), .Y(_4626_) );
NOR2X1 NOR2X1_69 ( .A(latched_rd_2_), .B(_4626_), .Y(_4627_) );
NAND2X1 NAND2X1_32 ( .A(_4624_), .B(_4627_), .Y(_4628_) );
INVX1 INVX1_66 ( .A(_4628_), .Y(_4629_) );
OAI21X1 OAI21X1_34 ( .A(latched_branch), .B(latched_store), .C(_4474_), .Y(_4630_) );
NOR2X1 NOR2X1_70 ( .A(_4630_), .B(_4629_), .Y(_4631_) );
INVX1 INVX1_67 ( .A(_4631_), .Y(_4632_) );
INVX1 INVX1_68 ( .A(latched_rd_3_), .Y(_4633_) );
NOR2X1 NOR2X1_71 ( .A(latched_rd_4_), .B(_4633_), .Y(_4634_) );
INVX1 INVX1_69 ( .A(_4634_), .Y(_4635_) );
NOR2X1 NOR2X1_72 ( .A(latched_rd_2_), .B(_4635_), .Y(_4636_) );
NAND2X1 NAND2X1_33 ( .A(_4624_), .B(_4636_), .Y(_4637_) );
NOR2X1 NOR2X1_73 ( .A(_4637__bF_buf3), .B(_4632__bF_buf8), .Y(_4638_) );
INVX1 INVX1_70 ( .A(latched_store), .Y(_4639_) );
NOR2X1 NOR2X1_74 ( .A(latched_branch), .B(_4639__bF_buf4), .Y(_4640_) );
INVX1 INVX1_71 ( .A(_4640_), .Y(_4641_) );
INVX1 INVX1_72 ( .A(reg_pc_4_), .Y(_4642_) );
INVX1 INVX1_73 ( .A(reg_pc_1_), .Y(_4643_) );
INVX1 INVX1_74 ( .A(reg_pc_2_), .Y(_4644_) );
AOI21X1 AOI21X1_7 ( .A(latched_compr), .B(_4643_), .C(_4644_), .Y(_4645_) );
NAND2X1 NAND2X1_34 ( .A(reg_pc_3_), .B(_4645_), .Y(_4646_) );
NOR2X1 NOR2X1_75 ( .A(_4642_), .B(_4646_), .Y(_4647_) );
NAND2X1 NAND2X1_35 ( .A(reg_pc_5_), .B(_4647_), .Y(_4648_) );
INVX1 INVX1_75 ( .A(_4648_), .Y(_4649_) );
NOR2X1 NOR2X1_76 ( .A(reg_pc_5_), .B(_4647_), .Y(_4650_) );
OAI21X1 OAI21X1_35 ( .A(_4649_), .B(_4650_), .C(_4641__bF_buf6), .Y(_4651_) );
MUX2X1 MUX2X1_2 ( .A(alu_out_q_5_), .B(reg_out_5_), .S(latched_stalu_bF_buf6), .Y(_4652_) );
INVX1 INVX1_76 ( .A(_4652_), .Y(_4653_) );
OAI21X1 OAI21X1_36 ( .A(_4641__bF_buf5), .B(_4653_), .C(_4651_), .Y(_4654_) );
INVX1 INVX1_77 ( .A(_4654__bF_buf4), .Y(_4655_) );
NAND2X1 NAND2X1_36 ( .A(_4638_), .B(_4655_), .Y(_4656_) );
OAI21X1 OAI21X1_37 ( .A(_4623_), .B(_4638_), .C(_4656_), .Y(_95_) );
INVX1 INVX1_78 ( .A(cpuregs_8_[6]), .Y(_4657_) );
INVX1 INVX1_79 ( .A(reg_pc_6_), .Y(_4658_) );
NOR2X1 NOR2X1_77 ( .A(_4658_), .B(_4648_), .Y(_4659_) );
NOR2X1 NOR2X1_78 ( .A(reg_pc_6_), .B(_4649_), .Y(_4660_) );
OAI21X1 OAI21X1_38 ( .A(_4660_), .B(_4659_), .C(_4641__bF_buf4), .Y(_4661_) );
MUX2X1 MUX2X1_3 ( .A(alu_out_q_6_), .B(reg_out_6_), .S(latched_stalu_bF_buf5), .Y(_4662_) );
INVX1 INVX1_80 ( .A(_4662_), .Y(_4663_) );
OAI21X1 OAI21X1_39 ( .A(_4641__bF_buf3), .B(_4663_), .C(_4661_), .Y(_4664_) );
INVX1 INVX1_81 ( .A(_4664__bF_buf4), .Y(_4665_) );
NAND2X1 NAND2X1_37 ( .A(_4638_), .B(_4665_), .Y(_4666_) );
OAI21X1 OAI21X1_40 ( .A(_4657_), .B(_4638_), .C(_4666_), .Y(_96_) );
INVX1 INVX1_82 ( .A(_4624_), .Y(_4667_) );
NAND2X1 NAND2X1_38 ( .A(_4636_), .B(_4631_), .Y(_4668_) );
NOR2X1 NOR2X1_79 ( .A(_4667_), .B(_4668_), .Y(_4669_) );
NOR2X1 NOR2X1_80 ( .A(cpuregs_8_[7]), .B(_4669_), .Y(_4670_) );
NAND2X1 NAND2X1_39 ( .A(reg_pc_7_), .B(_4659_), .Y(_4671_) );
INVX1 INVX1_83 ( .A(_4671_), .Y(_4672_) );
NOR2X1 NOR2X1_81 ( .A(reg_pc_7_), .B(_4659_), .Y(_4673_) );
OAI21X1 OAI21X1_41 ( .A(_4672_), .B(_4673_), .C(_4641__bF_buf2), .Y(_4674_) );
MUX2X1 MUX2X1_4 ( .A(alu_out_q_7_), .B(reg_out_7_), .S(latched_stalu_bF_buf4), .Y(_4675_) );
INVX1 INVX1_84 ( .A(_4675_), .Y(_4676_) );
OAI21X1 OAI21X1_42 ( .A(_4641__bF_buf1), .B(_4676_), .C(_4674_), .Y(_4677_) );
AOI21X1 AOI21X1_8 ( .A(_4669_), .B(_4677__bF_buf4), .C(_4670_), .Y(_97_) );
INVX1 INVX1_85 ( .A(cpuregs_8_[8]), .Y(_4678_) );
INVX1 INVX1_86 ( .A(reg_pc_8_), .Y(_4679_) );
NOR2X1 NOR2X1_82 ( .A(_4679_), .B(_4671_), .Y(_4680_) );
NOR2X1 NOR2X1_83 ( .A(reg_pc_8_), .B(_4672_), .Y(_4681_) );
OAI21X1 OAI21X1_43 ( .A(_4681_), .B(_4680_), .C(_4641__bF_buf0), .Y(_4682_) );
MUX2X1 MUX2X1_5 ( .A(alu_out_q_8_), .B(reg_out_8_), .S(latched_stalu_bF_buf3), .Y(_4683_) );
INVX1 INVX1_87 ( .A(_4683_), .Y(_4684_) );
OAI21X1 OAI21X1_44 ( .A(_4641__bF_buf6), .B(_4684_), .C(_4682_), .Y(_4685_) );
INVX1 INVX1_88 ( .A(_4685__bF_buf4), .Y(_4686_) );
NAND2X1 NAND2X1_40 ( .A(_4638_), .B(_4686_), .Y(_4687_) );
OAI21X1 OAI21X1_45 ( .A(_4678_), .B(_4638_), .C(_4687_), .Y(_98_) );
INVX1 INVX1_89 ( .A(cpuregs_8_[9]), .Y(_4688_) );
NAND2X1 NAND2X1_41 ( .A(reg_pc_8_), .B(reg_pc_9_), .Y(_4689_) );
NOR2X1 NOR2X1_84 ( .A(_4689_), .B(_4671_), .Y(_4690_) );
NOR2X1 NOR2X1_85 ( .A(reg_pc_9_), .B(_4680_), .Y(_4691_) );
OAI21X1 OAI21X1_46 ( .A(_4691_), .B(_4690_), .C(_4641__bF_buf5), .Y(_4692_) );
INVX1 INVX1_90 ( .A(reg_out_9_), .Y(_4693_) );
NAND2X1 NAND2X1_42 ( .A(latched_stalu_bF_buf2), .B(alu_out_q_9_), .Y(_4694_) );
OAI21X1 OAI21X1_47 ( .A(_4693_), .B(latched_stalu_bF_buf1), .C(_4694_), .Y(_4695_) );
OAI21X1 OAI21X1_48 ( .A(_4641__bF_buf4), .B(_4695_), .C(_4692_), .Y(_4696_) );
MUX2X1 MUX2X1_6 ( .A(_4696__bF_buf4), .B(_4688_), .S(_4669_), .Y(_99_) );
INVX1 INVX1_91 ( .A(cpuregs_8_[10]), .Y(_4697_) );
MUX2X1 MUX2X1_7 ( .A(alu_out_q_10_), .B(reg_out_10_), .S(latched_stalu_bF_buf0), .Y(_4698_) );
INVX1 INVX1_92 ( .A(_4698_), .Y(_4699_) );
NOR2X1 NOR2X1_86 ( .A(reg_pc_10_), .B(_4690_), .Y(_4700_) );
AND2X2 AND2X2_6 ( .A(_4690_), .B(reg_pc_10_), .Y(_4701_) );
OAI21X1 OAI21X1_49 ( .A(_4701_), .B(_4700_), .C(_4641__bF_buf3), .Y(_4702_) );
OAI21X1 OAI21X1_50 ( .A(_4641__bF_buf2), .B(_4699_), .C(_4702_), .Y(_4703_) );
MUX2X1 MUX2X1_8 ( .A(_4703__bF_buf4), .B(_4697_), .S(_4669_), .Y(_100_) );
INVX1 INVX1_93 ( .A(cpuregs_8_[11]), .Y(_4704_) );
MUX2X1 MUX2X1_9 ( .A(alu_out_q_11_), .B(reg_out_11_), .S(latched_stalu_bF_buf6), .Y(_4705_) );
INVX1 INVX1_94 ( .A(_4705_), .Y(_4706_) );
NOR2X1 NOR2X1_87 ( .A(reg_pc_11_), .B(_4701_), .Y(_4707_) );
NAND2X1 NAND2X1_43 ( .A(reg_pc_10_), .B(reg_pc_11_), .Y(_4708_) );
NOR2X1 NOR2X1_88 ( .A(_4689_), .B(_4708_), .Y(_4709_) );
NAND2X1 NAND2X1_44 ( .A(_4709_), .B(_4672_), .Y(_4710_) );
INVX1 INVX1_95 ( .A(_4710_), .Y(_4711_) );
OAI21X1 OAI21X1_51 ( .A(_4707_), .B(_4711_), .C(_4641__bF_buf1), .Y(_4712_) );
OAI21X1 OAI21X1_52 ( .A(_4641__bF_buf0), .B(_4706_), .C(_4712_), .Y(_4713_) );
MUX2X1 MUX2X1_10 ( .A(_4713__bF_buf4), .B(_4704_), .S(_4669_), .Y(_101_) );
INVX1 INVX1_96 ( .A(_4669_), .Y(_4714_) );
OAI21X1 OAI21X1_53 ( .A(_4632__bF_buf7), .B(_4637__bF_buf2), .C(cpuregs_8_[12]), .Y(_4715_) );
MUX2X1 MUX2X1_11 ( .A(alu_out_q_12_), .B(reg_out_12_), .S(latched_stalu_bF_buf5), .Y(_4716_) );
INVX1 INVX1_97 ( .A(_4716_), .Y(_4717_) );
NOR2X1 NOR2X1_89 ( .A(reg_pc_12_), .B(_4711_), .Y(_4718_) );
INVX1 INVX1_98 ( .A(reg_pc_12_), .Y(_4719_) );
NOR2X1 NOR2X1_90 ( .A(_4719_), .B(_4710_), .Y(_4720_) );
OAI21X1 OAI21X1_54 ( .A(_4718_), .B(_4720_), .C(_4641__bF_buf6), .Y(_4721_) );
OAI21X1 OAI21X1_55 ( .A(_4641__bF_buf5), .B(_4717_), .C(_4721_), .Y(_4722_) );
OAI21X1 OAI21X1_56 ( .A(_4722__bF_buf4), .B(_4714__bF_buf3), .C(_4715_), .Y(_102_) );
OAI21X1 OAI21X1_57 ( .A(_4632__bF_buf6), .B(_4637__bF_buf1), .C(cpuregs_8_[13]), .Y(_4723_) );
INVX1 INVX1_99 ( .A(reg_out_13_), .Y(_4724_) );
NAND2X1 NAND2X1_45 ( .A(latched_stalu_bF_buf4), .B(alu_out_q_13_), .Y(_4725_) );
OAI21X1 OAI21X1_58 ( .A(_4724_), .B(latched_stalu_bF_buf3), .C(_4725_), .Y(_4726_) );
NOR2X1 NOR2X1_91 ( .A(reg_pc_13_), .B(_4720_), .Y(_4727_) );
NAND2X1 NAND2X1_46 ( .A(reg_pc_13_), .B(_4720_), .Y(_4728_) );
INVX1 INVX1_100 ( .A(_4728_), .Y(_4729_) );
OAI21X1 OAI21X1_59 ( .A(_4729_), .B(_4727_), .C(_4641__bF_buf4), .Y(_4730_) );
OAI21X1 OAI21X1_60 ( .A(_4641__bF_buf3), .B(_4726_), .C(_4730_), .Y(_4731_) );
OAI21X1 OAI21X1_61 ( .A(_4731__bF_buf4), .B(_4714__bF_buf2), .C(_4723_), .Y(_103_) );
OAI21X1 OAI21X1_62 ( .A(_4632__bF_buf5), .B(_4637__bF_buf0), .C(cpuregs_8_[14]), .Y(_4732_) );
MUX2X1 MUX2X1_12 ( .A(alu_out_q_14_), .B(reg_out_14_), .S(latched_stalu_bF_buf2), .Y(_4733_) );
NAND2X1 NAND2X1_47 ( .A(_4733_), .B(_4640_), .Y(_4734_) );
NOR2X1 NOR2X1_92 ( .A(reg_pc_14_), .B(_4729_), .Y(_4735_) );
INVX1 INVX1_101 ( .A(reg_pc_14_), .Y(_4736_) );
NOR2X1 NOR2X1_93 ( .A(_4736_), .B(_4728_), .Y(_4737_) );
OAI21X1 OAI21X1_63 ( .A(_4735_), .B(_4737_), .C(_4641__bF_buf2), .Y(_4738_) );
AND2X2 AND2X2_7 ( .A(_4738_), .B(_4734_), .Y(_4739_) );
INVX1 INVX1_102 ( .A(_4739_), .Y(_4740_) );
OAI21X1 OAI21X1_64 ( .A(_4740__bF_buf4), .B(_4714__bF_buf1), .C(_4732_), .Y(_104_) );
OAI21X1 OAI21X1_65 ( .A(_4632__bF_buf4), .B(_4637__bF_buf3), .C(cpuregs_8_[15]), .Y(_4741_) );
MUX2X1 MUX2X1_13 ( .A(alu_out_q_15_), .B(reg_out_15_), .S(latched_stalu_bF_buf1), .Y(_4742_) );
INVX1 INVX1_103 ( .A(_4742_), .Y(_4743_) );
NOR2X1 NOR2X1_94 ( .A(reg_pc_15_), .B(_4737_), .Y(_4744_) );
AND2X2 AND2X2_8 ( .A(_4737_), .B(reg_pc_15_), .Y(_4745_) );
OAI21X1 OAI21X1_66 ( .A(_4745_), .B(_4744_), .C(_4641__bF_buf1), .Y(_4746_) );
OAI21X1 OAI21X1_67 ( .A(_4641__bF_buf0), .B(_4743_), .C(_4746_), .Y(_4747_) );
OAI21X1 OAI21X1_68 ( .A(_4747__bF_buf4), .B(_4714__bF_buf0), .C(_4741_), .Y(_105_) );
OAI21X1 OAI21X1_69 ( .A(_4632__bF_buf3), .B(_4637__bF_buf2), .C(cpuregs_8_[16]), .Y(_4748_) );
INVX1 INVX1_104 ( .A(reg_out_16_), .Y(_4749_) );
NAND2X1 NAND2X1_48 ( .A(latched_stalu_bF_buf0), .B(alu_out_q_16_), .Y(_4750_) );
OAI21X1 OAI21X1_70 ( .A(_4749_), .B(latched_stalu_bF_buf6), .C(_4750_), .Y(_4751_) );
NOR2X1 NOR2X1_95 ( .A(reg_pc_16_), .B(_4745_), .Y(_4752_) );
AND2X2 AND2X2_9 ( .A(_4745_), .B(reg_pc_16_), .Y(_4753_) );
OAI21X1 OAI21X1_71 ( .A(_4753_), .B(_4752_), .C(_4641__bF_buf6), .Y(_4754_) );
OAI21X1 OAI21X1_72 ( .A(_4641__bF_buf5), .B(_4751_), .C(_4754_), .Y(_4755_) );
OAI21X1 OAI21X1_73 ( .A(_4755__bF_buf4), .B(_4714__bF_buf3), .C(_4748_), .Y(_106_) );
OAI21X1 OAI21X1_74 ( .A(_4632__bF_buf2), .B(_4637__bF_buf1), .C(cpuregs_8_[17]), .Y(_4756_) );
INVX1 INVX1_105 ( .A(reg_out_17_), .Y(_4757_) );
NAND2X1 NAND2X1_49 ( .A(latched_stalu_bF_buf5), .B(alu_out_q_17_), .Y(_4758_) );
OAI21X1 OAI21X1_75 ( .A(_4757_), .B(latched_stalu_bF_buf4), .C(_4758_), .Y(_4759_) );
NOR2X1 NOR2X1_96 ( .A(reg_pc_17_), .B(_4753_), .Y(_4760_) );
AND2X2 AND2X2_10 ( .A(_4753_), .B(reg_pc_17_), .Y(_4761_) );
OAI21X1 OAI21X1_76 ( .A(_4761_), .B(_4760_), .C(_4641__bF_buf4), .Y(_4762_) );
OAI21X1 OAI21X1_77 ( .A(_4641__bF_buf3), .B(_4759_), .C(_4762_), .Y(_4763_) );
OAI21X1 OAI21X1_78 ( .A(_4763__bF_buf4), .B(_4714__bF_buf2), .C(_4756_), .Y(_107_) );
OAI21X1 OAI21X1_79 ( .A(_4632__bF_buf1), .B(_4637__bF_buf0), .C(cpuregs_8_[18]), .Y(_4764_) );
INVX1 INVX1_106 ( .A(reg_out_18_), .Y(_4765_) );
NAND2X1 NAND2X1_50 ( .A(latched_stalu_bF_buf3), .B(alu_out_q_18_), .Y(_4766_) );
OAI21X1 OAI21X1_80 ( .A(_4765_), .B(latched_stalu_bF_buf2), .C(_4766_), .Y(_4767_) );
INVX1 INVX1_107 ( .A(reg_pc_13_), .Y(_4768_) );
NOR2X1 NOR2X1_97 ( .A(_4719_), .B(_4768_), .Y(_4769_) );
AND2X2 AND2X2_11 ( .A(reg_pc_14_), .B(reg_pc_15_), .Y(_4770_) );
NAND3X1 NAND3X1_10 ( .A(_4769_), .B(_4770_), .C(_4709_), .Y(_4771_) );
NOR2X1 NOR2X1_98 ( .A(_4771_), .B(_4671_), .Y(_4772_) );
INVX1 INVX1_108 ( .A(_4772_), .Y(_4773_) );
INVX1 INVX1_109 ( .A(reg_pc_16_), .Y(_4774_) );
INVX1 INVX1_110 ( .A(reg_pc_17_), .Y(_4775_) );
NOR2X1 NOR2X1_99 ( .A(_4774_), .B(_4775_), .Y(_4776_) );
INVX1 INVX1_111 ( .A(_4776_), .Y(_4777_) );
OAI21X1 OAI21X1_81 ( .A(_4773_), .B(_4777_), .C(reg_pc_18_), .Y(_4778_) );
INVX1 INVX1_112 ( .A(reg_pc_18_), .Y(_4779_) );
NOR2X1 NOR2X1_100 ( .A(_4777_), .B(_4773_), .Y(_4780_) );
NAND2X1 NAND2X1_51 ( .A(_4779_), .B(_4780_), .Y(_4781_) );
NAND3X1 NAND3X1_11 ( .A(_4641__bF_buf2), .B(_4778_), .C(_4781_), .Y(_4782_) );
OAI21X1 OAI21X1_82 ( .A(_4641__bF_buf1), .B(_4767_), .C(_4782_), .Y(_4783_) );
OAI21X1 OAI21X1_83 ( .A(_4783__bF_buf4), .B(_4714__bF_buf1), .C(_4764_), .Y(_108_) );
OAI21X1 OAI21X1_84 ( .A(_4632__bF_buf0), .B(_4637__bF_buf3), .C(cpuregs_8_[19]), .Y(_4784_) );
INVX1 INVX1_113 ( .A(reg_out_19_), .Y(_4785_) );
NAND2X1 NAND2X1_52 ( .A(latched_stalu_bF_buf1), .B(alu_out_q_19_), .Y(_4786_) );
OAI21X1 OAI21X1_85 ( .A(_4785_), .B(latched_stalu_bF_buf0), .C(_4786_), .Y(_4787_) );
INVX1 INVX1_114 ( .A(_4780_), .Y(_4788_) );
OAI21X1 OAI21X1_86 ( .A(_4788_), .B(_4779_), .C(reg_pc_19_), .Y(_4789_) );
INVX1 INVX1_115 ( .A(reg_pc_19_), .Y(_4790_) );
NAND3X1 NAND3X1_12 ( .A(reg_pc_18_), .B(_4790_), .C(_4780_), .Y(_4791_) );
NAND3X1 NAND3X1_13 ( .A(_4641__bF_buf0), .B(_4791_), .C(_4789_), .Y(_4792_) );
OAI21X1 OAI21X1_87 ( .A(_4641__bF_buf6), .B(_4787_), .C(_4792_), .Y(_4793_) );
OAI21X1 OAI21X1_88 ( .A(_4793__bF_buf4), .B(_4714__bF_buf0), .C(_4784_), .Y(_109_) );
OAI21X1 OAI21X1_89 ( .A(_4632__bF_buf8), .B(_4637__bF_buf2), .C(cpuregs_8_[20]), .Y(_4794_) );
INVX1 INVX1_116 ( .A(reg_out_20_), .Y(_4795_) );
NAND2X1 NAND2X1_53 ( .A(latched_stalu_bF_buf6), .B(alu_out_q_20_), .Y(_4796_) );
OAI21X1 OAI21X1_90 ( .A(_4795_), .B(latched_stalu_bF_buf5), .C(_4796_), .Y(_4797_) );
NAND2X1 NAND2X1_54 ( .A(reg_pc_18_), .B(reg_pc_19_), .Y(_4798_) );
NOR2X1 NOR2X1_101 ( .A(_4798_), .B(_4777_), .Y(_4799_) );
NAND2X1 NAND2X1_55 ( .A(_4799_), .B(_4772_), .Y(_4800_) );
INVX1 INVX1_117 ( .A(_4800_), .Y(_4801_) );
NOR2X1 NOR2X1_102 ( .A(reg_pc_20_), .B(_4801_), .Y(_4802_) );
INVX1 INVX1_118 ( .A(reg_pc_20_), .Y(_4803_) );
NOR2X1 NOR2X1_103 ( .A(_4803_), .B(_4800_), .Y(_4804_) );
OAI21X1 OAI21X1_91 ( .A(_4802_), .B(_4804_), .C(_4641__bF_buf5), .Y(_4805_) );
OAI21X1 OAI21X1_92 ( .A(_4641__bF_buf4), .B(_4797_), .C(_4805_), .Y(_4806_) );
OAI21X1 OAI21X1_93 ( .A(_4806__bF_buf4), .B(_4714__bF_buf3), .C(_4794_), .Y(_110_) );
OAI21X1 OAI21X1_94 ( .A(_4632__bF_buf7), .B(_4637__bF_buf1), .C(cpuregs_8_[21]), .Y(_4807_) );
INVX1 INVX1_119 ( .A(reg_out_21_), .Y(_4808_) );
NAND2X1 NAND2X1_56 ( .A(latched_stalu_bF_buf4), .B(alu_out_q_21_), .Y(_4809_) );
OAI21X1 OAI21X1_95 ( .A(_4808_), .B(latched_stalu_bF_buf3), .C(_4809_), .Y(_4810_) );
NOR2X1 NOR2X1_104 ( .A(reg_pc_21_), .B(_4804_), .Y(_4811_) );
INVX1 INVX1_120 ( .A(reg_pc_21_), .Y(_4812_) );
INVX1 INVX1_121 ( .A(_4804_), .Y(_4813_) );
NOR2X1 NOR2X1_105 ( .A(_4812_), .B(_4813_), .Y(_4814_) );
OAI21X1 OAI21X1_96 ( .A(_4814_), .B(_4811_), .C(_4641__bF_buf3), .Y(_4815_) );
OAI21X1 OAI21X1_97 ( .A(_4641__bF_buf2), .B(_4810_), .C(_4815_), .Y(_4816_) );
OAI21X1 OAI21X1_98 ( .A(_4816__bF_buf4), .B(_4714__bF_buf2), .C(_4807_), .Y(_111_) );
OAI21X1 OAI21X1_99 ( .A(_4632__bF_buf6), .B(_4637__bF_buf0), .C(cpuregs_8_[22]), .Y(_4817_) );
INVX1 INVX1_122 ( .A(reg_out_22_), .Y(_4818_) );
NAND2X1 NAND2X1_57 ( .A(latched_stalu_bF_buf2), .B(alu_out_q_22_), .Y(_4819_) );
OAI21X1 OAI21X1_100 ( .A(_4818_), .B(latched_stalu_bF_buf1), .C(_4819_), .Y(_4820_) );
NOR2X1 NOR2X1_106 ( .A(reg_pc_22_), .B(_4814_), .Y(_4821_) );
AND2X2 AND2X2_12 ( .A(_4814_), .B(reg_pc_22_), .Y(_4822_) );
OAI21X1 OAI21X1_101 ( .A(_4822_), .B(_4821_), .C(_4641__bF_buf1), .Y(_4823_) );
OAI21X1 OAI21X1_102 ( .A(_4641__bF_buf0), .B(_4820_), .C(_4823_), .Y(_4824_) );
OAI21X1 OAI21X1_103 ( .A(_4824__bF_buf4), .B(_4714__bF_buf1), .C(_4817_), .Y(_112_) );
OAI21X1 OAI21X1_104 ( .A(_4632__bF_buf5), .B(_4637__bF_buf3), .C(cpuregs_8_[23]), .Y(_4825_) );
INVX1 INVX1_123 ( .A(reg_pc_23_), .Y(_4826_) );
XNOR2X1 XNOR2X1_1 ( .A(_4822_), .B(_4826_), .Y(_4827_) );
INVX1 INVX1_124 ( .A(reg_out_23_), .Y(_4828_) );
NAND2X1 NAND2X1_58 ( .A(latched_stalu_bF_buf0), .B(alu_out_q_23_), .Y(_4829_) );
OAI21X1 OAI21X1_105 ( .A(_4828_), .B(latched_stalu_bF_buf6), .C(_4829_), .Y(_4830_) );
INVX1 INVX1_125 ( .A(_4830_), .Y(_4831_) );
NAND2X1 NAND2X1_59 ( .A(_4640_), .B(_4831_), .Y(_4832_) );
OAI21X1 OAI21X1_106 ( .A(_4827_), .B(_4640_), .C(_4832_), .Y(_4833_) );
OAI21X1 OAI21X1_107 ( .A(_4833__bF_buf4), .B(_4714__bF_buf0), .C(_4825_), .Y(_113_) );
OAI21X1 OAI21X1_108 ( .A(_4632__bF_buf4), .B(_4637__bF_buf2), .C(cpuregs_8_[24]), .Y(_4834_) );
INVX1 INVX1_126 ( .A(reg_out_24_), .Y(_4835_) );
NAND2X1 NAND2X1_60 ( .A(latched_stalu_bF_buf5), .B(alu_out_q_24_), .Y(_4836_) );
OAI21X1 OAI21X1_109 ( .A(_4835_), .B(latched_stalu_bF_buf4), .C(_4836_), .Y(_4837_) );
NAND3X1 NAND3X1_14 ( .A(reg_pc_21_), .B(reg_pc_22_), .C(reg_pc_23_), .Y(_4838_) );
INVX1 INVX1_127 ( .A(_4838_), .Y(_4839_) );
AOI21X1 AOI21X1_9 ( .A(_4839_), .B(_4804_), .C(reg_pc_24_), .Y(_4840_) );
INVX1 INVX1_128 ( .A(reg_pc_24_), .Y(_4841_) );
NAND2X1 NAND2X1_61 ( .A(_4839_), .B(_4804_), .Y(_4842_) );
NOR2X1 NOR2X1_107 ( .A(_4841_), .B(_4842_), .Y(_4843_) );
OAI21X1 OAI21X1_110 ( .A(_4843_), .B(_4840_), .C(_4641__bF_buf6), .Y(_4844_) );
OAI21X1 OAI21X1_111 ( .A(_4641__bF_buf5), .B(_4837_), .C(_4844_), .Y(_4845_) );
OAI21X1 OAI21X1_112 ( .A(_4845__bF_buf4), .B(_4714__bF_buf3), .C(_4834_), .Y(_114_) );
OAI21X1 OAI21X1_113 ( .A(_4632__bF_buf3), .B(_4637__bF_buf1), .C(cpuregs_8_[25]), .Y(_4846_) );
INVX1 INVX1_129 ( .A(reg_out_25_), .Y(_4847_) );
NAND2X1 NAND2X1_62 ( .A(latched_stalu_bF_buf3), .B(alu_out_q_25_), .Y(_4848_) );
OAI21X1 OAI21X1_114 ( .A(_4847_), .B(latched_stalu_bF_buf2), .C(_4848_), .Y(_4849_) );
NOR2X1 NOR2X1_108 ( .A(reg_pc_25_), .B(_4843_), .Y(_4850_) );
NAND2X1 NAND2X1_63 ( .A(reg_pc_25_), .B(_4843_), .Y(_4851_) );
INVX1 INVX1_130 ( .A(_4851_), .Y(_4852_) );
OAI21X1 OAI21X1_115 ( .A(_4852_), .B(_4850_), .C(_4641__bF_buf4), .Y(_4853_) );
OAI21X1 OAI21X1_116 ( .A(_4641__bF_buf3), .B(_4849_), .C(_4853_), .Y(_4854_) );
OAI21X1 OAI21X1_117 ( .A(_4854__bF_buf4), .B(_4714__bF_buf2), .C(_4846_), .Y(_115_) );
OAI21X1 OAI21X1_118 ( .A(_4632__bF_buf2), .B(_4637__bF_buf0), .C(cpuregs_8_[26]), .Y(_4855_) );
INVX1 INVX1_131 ( .A(reg_out_26_), .Y(_4856_) );
NAND2X1 NAND2X1_64 ( .A(latched_stalu_bF_buf1), .B(alu_out_q_26_), .Y(_4857_) );
OAI21X1 OAI21X1_119 ( .A(_4856_), .B(latched_stalu_bF_buf0), .C(_4857_), .Y(_4858_) );
NOR2X1 NOR2X1_109 ( .A(reg_pc_26_), .B(_4852_), .Y(_4859_) );
INVX1 INVX1_132 ( .A(reg_pc_26_), .Y(_4860_) );
NOR2X1 NOR2X1_110 ( .A(_4860_), .B(_4851_), .Y(_4861_) );
OAI21X1 OAI21X1_120 ( .A(_4859_), .B(_4861_), .C(_4641__bF_buf2), .Y(_4862_) );
OAI21X1 OAI21X1_121 ( .A(_4641__bF_buf1), .B(_4858_), .C(_4862_), .Y(_4863_) );
OAI21X1 OAI21X1_122 ( .A(_4863__bF_buf4), .B(_4714__bF_buf1), .C(_4855_), .Y(_116_) );
OAI21X1 OAI21X1_123 ( .A(_4632__bF_buf1), .B(_4637__bF_buf3), .C(cpuregs_8_[27]), .Y(_4864_) );
XOR2X1 XOR2X1_1 ( .A(_4861_), .B(reg_pc_27_), .Y(_4865_) );
INVX1 INVX1_133 ( .A(reg_out_27_), .Y(_4866_) );
NAND2X1 NAND2X1_65 ( .A(latched_stalu_bF_buf6), .B(alu_out_q_27_), .Y(_4867_) );
OAI21X1 OAI21X1_124 ( .A(_4866_), .B(latched_stalu_bF_buf5), .C(_4867_), .Y(_4868_) );
INVX1 INVX1_134 ( .A(_4868_), .Y(_4869_) );
NAND2X1 NAND2X1_66 ( .A(_4640_), .B(_4869_), .Y(_4870_) );
OAI21X1 OAI21X1_125 ( .A(_4865_), .B(_4640_), .C(_4870_), .Y(_4871_) );
OAI21X1 OAI21X1_126 ( .A(_4871__bF_buf4), .B(_4714__bF_buf0), .C(_4864_), .Y(_117_) );
OAI21X1 OAI21X1_127 ( .A(_4632__bF_buf0), .B(_4637__bF_buf2), .C(cpuregs_8_[28]), .Y(_4872_) );
INVX1 INVX1_135 ( .A(reg_out_28_), .Y(_4873_) );
NAND2X1 NAND2X1_67 ( .A(latched_stalu_bF_buf4), .B(alu_out_q_28_), .Y(_4874_) );
OAI21X1 OAI21X1_128 ( .A(_4873_), .B(latched_stalu_bF_buf3), .C(_4874_), .Y(_4875_) );
AOI21X1 AOI21X1_10 ( .A(reg_pc_27_), .B(_4861_), .C(reg_pc_28_), .Y(_4876_) );
INVX1 INVX1_136 ( .A(reg_pc_25_), .Y(_4877_) );
NOR2X1 NOR2X1_111 ( .A(_4841_), .B(_4877_), .Y(_4878_) );
NAND3X1 NAND3X1_15 ( .A(reg_pc_26_), .B(reg_pc_27_), .C(_4878_), .Y(_4879_) );
NOR2X1 NOR2X1_112 ( .A(_4879_), .B(_4842_), .Y(_4880_) );
NAND2X1 NAND2X1_68 ( .A(reg_pc_28_), .B(_4880_), .Y(_4881_) );
INVX1 INVX1_137 ( .A(_4881_), .Y(_4882_) );
OAI21X1 OAI21X1_129 ( .A(_4876_), .B(_4882_), .C(_4641__bF_buf0), .Y(_4883_) );
OAI21X1 OAI21X1_130 ( .A(_4641__bF_buf6), .B(_4875_), .C(_4883_), .Y(_4884_) );
OAI21X1 OAI21X1_131 ( .A(_4884__bF_buf4), .B(_4714__bF_buf3), .C(_4872_), .Y(_118_) );
OAI21X1 OAI21X1_132 ( .A(_4632__bF_buf8), .B(_4637__bF_buf1), .C(cpuregs_8_[29]), .Y(_4885_) );
INVX1 INVX1_138 ( .A(reg_out_29_), .Y(_4886_) );
NAND2X1 NAND2X1_69 ( .A(latched_stalu_bF_buf2), .B(alu_out_q_29_), .Y(_4887_) );
OAI21X1 OAI21X1_133 ( .A(_4886_), .B(latched_stalu_bF_buf1), .C(_4887_), .Y(_4888_) );
NOR2X1 NOR2X1_113 ( .A(reg_pc_29_), .B(_4882_), .Y(_4889_) );
INVX1 INVX1_139 ( .A(reg_pc_29_), .Y(_4890_) );
NOR2X1 NOR2X1_114 ( .A(_4890_), .B(_4881_), .Y(_4891_) );
OAI21X1 OAI21X1_134 ( .A(_4889_), .B(_4891_), .C(_4641__bF_buf5), .Y(_4892_) );
OAI21X1 OAI21X1_135 ( .A(_4641__bF_buf4), .B(_4888_), .C(_4892_), .Y(_4893_) );
OAI21X1 OAI21X1_136 ( .A(_4893__bF_buf4), .B(_4714__bF_buf2), .C(_4885_), .Y(_119_) );
OAI21X1 OAI21X1_137 ( .A(_4632__bF_buf7), .B(_4637__bF_buf0), .C(cpuregs_8_[30]), .Y(_4894_) );
INVX1 INVX1_140 ( .A(reg_out_30_), .Y(_4895_) );
NAND2X1 NAND2X1_70 ( .A(latched_stalu_bF_buf0), .B(alu_out_q_30_), .Y(_4896_) );
OAI21X1 OAI21X1_138 ( .A(_4895_), .B(latched_stalu_bF_buf6), .C(_4896_), .Y(_4897_) );
INVX1 INVX1_141 ( .A(reg_pc_30_), .Y(_4898_) );
OAI21X1 OAI21X1_139 ( .A(_4881_), .B(_4890_), .C(_4898_), .Y(_4899_) );
AOI21X1 AOI21X1_11 ( .A(reg_pc_30_), .B(_4891_), .C(_4640_), .Y(_4900_) );
AOI22X1 AOI22X1_4 ( .A(_4640_), .B(_4897_), .C(_4900_), .D(_4899_), .Y(_4901_) );
OAI21X1 OAI21X1_140 ( .A(_4901__bF_buf4), .B(_4714__bF_buf1), .C(_4894_), .Y(_120_) );
OAI21X1 OAI21X1_141 ( .A(_4632__bF_buf6), .B(_4637__bF_buf3), .C(cpuregs_8_[31]), .Y(_4902_) );
INVX1 INVX1_142 ( .A(reg_out_31_), .Y(_4903_) );
NAND2X1 NAND2X1_71 ( .A(latched_stalu_bF_buf5), .B(alu_out_q_31_), .Y(_4904_) );
OAI21X1 OAI21X1_142 ( .A(_4903_), .B(latched_stalu_bF_buf4), .C(_4904_), .Y(_4905_) );
NAND3X1 NAND3X1_16 ( .A(reg_pc_30_), .B(reg_pc_31_), .C(_4891_), .Y(_4906_) );
INVX1 INVX1_143 ( .A(reg_pc_31_), .Y(_4907_) );
NAND2X1 NAND2X1_72 ( .A(reg_pc_30_), .B(_4891_), .Y(_4908_) );
AOI21X1 AOI21X1_12 ( .A(_4907_), .B(_4908_), .C(_4640_), .Y(_4909_) );
AOI22X1 AOI22X1_5 ( .A(_4640_), .B(_4905_), .C(_4909_), .D(_4906_), .Y(_4910_) );
OAI21X1 OAI21X1_143 ( .A(_4910__bF_buf4), .B(_4714__bF_buf0), .C(_4902_), .Y(_121_) );
INVX1 INVX1_144 ( .A(latched_rd_2_), .Y(_4911_) );
NOR2X1 NOR2X1_115 ( .A(_4911_), .B(_4626_), .Y(_4912_) );
INVX1 INVX1_145 ( .A(_4912_), .Y(_4913_) );
INVX1 INVX1_146 ( .A(latched_rd_1_), .Y(_4914_) );
INVX1 INVX1_147 ( .A(latched_rd_0_), .Y(_4915_) );
NOR2X1 NOR2X1_116 ( .A(_4914_), .B(_4915_), .Y(_4916_) );
NAND2X1 NAND2X1_73 ( .A(_4916_), .B(_4631_), .Y(_4917_) );
NOR2X1 NOR2X1_117 ( .A(_4913__bF_buf6), .B(_4917__bF_buf10), .Y(_4918_) );
INVX1 INVX1_148 ( .A(_4918_), .Y(_4919_) );
INVX1 INVX1_149 ( .A(reg_out_0_), .Y(_4920_) );
NAND2X1 NAND2X1_74 ( .A(latched_stalu_bF_buf3), .B(alu_out_q_0_), .Y(_4921_) );
OAI21X1 OAI21X1_144 ( .A(_4920_), .B(latched_stalu_bF_buf2), .C(_4921_), .Y(_4922_) );
INVX1 INVX1_150 ( .A(reg_pc_0_), .Y(_4923_) );
OAI21X1 OAI21X1_145 ( .A(_4639__bF_buf3), .B(latched_branch), .C(_4923_), .Y(_4924_) );
OAI21X1 OAI21X1_146 ( .A(_4641__bF_buf3), .B(_4922_), .C(_4924_), .Y(_4925_) );
OAI21X1 OAI21X1_147 ( .A(_4917__bF_buf9), .B(_4913__bF_buf5), .C(cpuregs_7_[0]), .Y(_4926_) );
OAI21X1 OAI21X1_148 ( .A(_4919__bF_buf4), .B(_4925__bF_buf4), .C(_4926_), .Y(_122_) );
NOR2X1 NOR2X1_118 ( .A(latched_compr), .B(_4643_), .Y(_4927_) );
NAND2X1 NAND2X1_75 ( .A(latched_compr), .B(_4643_), .Y(_4928_) );
OAI21X1 OAI21X1_149 ( .A(latched_branch), .B(_4639__bF_buf2), .C(_4928_), .Y(_4929_) );
INVX1 INVX1_151 ( .A(reg_out_1_), .Y(_4930_) );
NAND2X1 NAND2X1_76 ( .A(latched_stalu_bF_buf1), .B(alu_out_q_1_), .Y(_4931_) );
OAI21X1 OAI21X1_150 ( .A(_4930_), .B(latched_stalu_bF_buf0), .C(_4931_), .Y(_4932_) );
OAI22X1 OAI22X1_3 ( .A(_4641__bF_buf2), .B(_4932_), .C(_4929_), .D(_4927_), .Y(_4933_) );
OAI21X1 OAI21X1_151 ( .A(_4917__bF_buf8), .B(_4913__bF_buf4), .C(cpuregs_7_[1]), .Y(_4934_) );
OAI21X1 OAI21X1_152 ( .A(_4919__bF_buf3), .B(_4933__bF_buf4), .C(_4934_), .Y(_123_) );
NOR2X1 NOR2X1_119 ( .A(reg_pc_2_), .B(_4928_), .Y(_4935_) );
OAI21X1 OAI21X1_153 ( .A(_4935_), .B(_4645_), .C(_4641__bF_buf1), .Y(_4936_) );
INVX1 INVX1_152 ( .A(reg_out_2_), .Y(_4937_) );
NAND2X1 NAND2X1_77 ( .A(latched_stalu_bF_buf6), .B(alu_out_q_2_), .Y(_4938_) );
OAI21X1 OAI21X1_154 ( .A(_4937_), .B(latched_stalu_bF_buf5), .C(_4938_), .Y(_4939_) );
OAI21X1 OAI21X1_155 ( .A(_4641__bF_buf0), .B(_4939_), .C(_4936_), .Y(_4940_) );
OAI21X1 OAI21X1_156 ( .A(_4917__bF_buf7), .B(_4913__bF_buf3), .C(cpuregs_7_[2]), .Y(_4941_) );
OAI21X1 OAI21X1_157 ( .A(_4919__bF_buf2), .B(_4940__bF_buf4), .C(_4941_), .Y(_124_) );
INVX1 INVX1_153 ( .A(_4646_), .Y(_4942_) );
NOR2X1 NOR2X1_120 ( .A(reg_pc_3_), .B(_4645_), .Y(_4943_) );
OAI21X1 OAI21X1_158 ( .A(_4942_), .B(_4943_), .C(_4641__bF_buf6), .Y(_4944_) );
INVX1 INVX1_154 ( .A(reg_out_3_), .Y(_4945_) );
NAND2X1 NAND2X1_78 ( .A(latched_stalu_bF_buf4), .B(alu_out_q_3_), .Y(_4946_) );
OAI21X1 OAI21X1_159 ( .A(_4945_), .B(latched_stalu_bF_buf3), .C(_4946_), .Y(_4947_) );
OAI21X1 OAI21X1_160 ( .A(_4641__bF_buf5), .B(_4947_), .C(_4944_), .Y(_4948_) );
OAI21X1 OAI21X1_161 ( .A(_4917__bF_buf6), .B(_4913__bF_buf2), .C(cpuregs_7_[3]), .Y(_4949_) );
OAI21X1 OAI21X1_162 ( .A(_4919__bF_buf1), .B(_4948__bF_buf4), .C(_4949_), .Y(_125_) );
NOR2X1 NOR2X1_121 ( .A(reg_pc_4_), .B(_4942_), .Y(_4950_) );
OAI21X1 OAI21X1_163 ( .A(_4950_), .B(_4647_), .C(_4641__bF_buf4), .Y(_4951_) );
INVX1 INVX1_155 ( .A(reg_out_4_), .Y(_4952_) );
NAND2X1 NAND2X1_79 ( .A(latched_stalu_bF_buf2), .B(alu_out_q_4_), .Y(_4953_) );
OAI21X1 OAI21X1_164 ( .A(_4952_), .B(latched_stalu_bF_buf1), .C(_4953_), .Y(_4954_) );
OAI21X1 OAI21X1_165 ( .A(_4641__bF_buf3), .B(_4954_), .C(_4951_), .Y(_4955_) );
OAI21X1 OAI21X1_166 ( .A(_4917__bF_buf5), .B(_4913__bF_buf1), .C(cpuregs_7_[4]), .Y(_4956_) );
OAI21X1 OAI21X1_167 ( .A(_4919__bF_buf0), .B(_4955__bF_buf4), .C(_4956_), .Y(_126_) );
OAI21X1 OAI21X1_168 ( .A(_4917__bF_buf4), .B(_4913__bF_buf0), .C(cpuregs_7_[5]), .Y(_4957_) );
OAI21X1 OAI21X1_169 ( .A(_4919__bF_buf4), .B(_4654__bF_buf3), .C(_4957_), .Y(_127_) );
OAI21X1 OAI21X1_170 ( .A(_4917__bF_buf3), .B(_4913__bF_buf6), .C(cpuregs_7_[6]), .Y(_4958_) );
OAI21X1 OAI21X1_171 ( .A(_4664__bF_buf3), .B(_4919__bF_buf3), .C(_4958_), .Y(_128_) );
OAI21X1 OAI21X1_172 ( .A(_4917__bF_buf2), .B(_4913__bF_buf5), .C(cpuregs_7_[7]), .Y(_4959_) );
OAI21X1 OAI21X1_173 ( .A(_4677__bF_buf3), .B(_4919__bF_buf2), .C(_4959_), .Y(_129_) );
OAI21X1 OAI21X1_174 ( .A(_4917__bF_buf1), .B(_4913__bF_buf4), .C(cpuregs_7_[8]), .Y(_4960_) );
OAI21X1 OAI21X1_175 ( .A(_4685__bF_buf3), .B(_4919__bF_buf1), .C(_4960_), .Y(_130_) );
OAI21X1 OAI21X1_176 ( .A(_4917__bF_buf0), .B(_4913__bF_buf3), .C(cpuregs_7_[9]), .Y(_4961_) );
OAI21X1 OAI21X1_177 ( .A(_4696__bF_buf3), .B(_4919__bF_buf0), .C(_4961_), .Y(_131_) );
OAI21X1 OAI21X1_178 ( .A(_4917__bF_buf10), .B(_4913__bF_buf2), .C(cpuregs_7_[10]), .Y(_4962_) );
OAI21X1 OAI21X1_179 ( .A(_4703__bF_buf3), .B(_4919__bF_buf4), .C(_4962_), .Y(_132_) );
OAI21X1 OAI21X1_180 ( .A(_4917__bF_buf9), .B(_4913__bF_buf1), .C(cpuregs_7_[11]), .Y(_4963_) );
OAI21X1 OAI21X1_181 ( .A(_4713__bF_buf3), .B(_4919__bF_buf3), .C(_4963_), .Y(_133_) );
OAI21X1 OAI21X1_182 ( .A(_4917__bF_buf8), .B(_4913__bF_buf0), .C(cpuregs_7_[12]), .Y(_4964_) );
OAI21X1 OAI21X1_183 ( .A(_4722__bF_buf3), .B(_4919__bF_buf2), .C(_4964_), .Y(_134_) );
OAI21X1 OAI21X1_184 ( .A(_4917__bF_buf7), .B(_4913__bF_buf6), .C(cpuregs_7_[13]), .Y(_4965_) );
OAI21X1 OAI21X1_185 ( .A(_4731__bF_buf3), .B(_4919__bF_buf1), .C(_4965_), .Y(_135_) );
OAI21X1 OAI21X1_186 ( .A(_4917__bF_buf6), .B(_4913__bF_buf5), .C(cpuregs_7_[14]), .Y(_4966_) );
OAI21X1 OAI21X1_187 ( .A(_4740__bF_buf3), .B(_4919__bF_buf0), .C(_4966_), .Y(_136_) );
OAI21X1 OAI21X1_188 ( .A(_4917__bF_buf5), .B(_4913__bF_buf4), .C(cpuregs_7_[15]), .Y(_4967_) );
OAI21X1 OAI21X1_189 ( .A(_4747__bF_buf3), .B(_4919__bF_buf4), .C(_4967_), .Y(_137_) );
OAI21X1 OAI21X1_190 ( .A(_4917__bF_buf4), .B(_4913__bF_buf3), .C(cpuregs_7_[16]), .Y(_4968_) );
OAI21X1 OAI21X1_191 ( .A(_4755__bF_buf3), .B(_4919__bF_buf3), .C(_4968_), .Y(_138_) );
OAI21X1 OAI21X1_192 ( .A(_4917__bF_buf3), .B(_4913__bF_buf2), .C(cpuregs_7_[17]), .Y(_4969_) );
OAI21X1 OAI21X1_193 ( .A(_4763__bF_buf3), .B(_4919__bF_buf2), .C(_4969_), .Y(_139_) );
OAI21X1 OAI21X1_194 ( .A(_4917__bF_buf2), .B(_4913__bF_buf1), .C(cpuregs_7_[18]), .Y(_4970_) );
OAI21X1 OAI21X1_195 ( .A(_4783__bF_buf3), .B(_4919__bF_buf1), .C(_4970_), .Y(_140_) );
OAI21X1 OAI21X1_196 ( .A(_4917__bF_buf1), .B(_4913__bF_buf0), .C(cpuregs_7_[19]), .Y(_4971_) );
OAI21X1 OAI21X1_197 ( .A(_4793__bF_buf3), .B(_4919__bF_buf0), .C(_4971_), .Y(_141_) );
OAI21X1 OAI21X1_198 ( .A(_4917__bF_buf0), .B(_4913__bF_buf6), .C(cpuregs_7_[20]), .Y(_4972_) );
OAI21X1 OAI21X1_199 ( .A(_4806__bF_buf3), .B(_4919__bF_buf4), .C(_4972_), .Y(_142_) );
OAI21X1 OAI21X1_200 ( .A(_4917__bF_buf10), .B(_4913__bF_buf5), .C(cpuregs_7_[21]), .Y(_4973_) );
OAI21X1 OAI21X1_201 ( .A(_4816__bF_buf3), .B(_4919__bF_buf3), .C(_4973_), .Y(_143_) );
OAI21X1 OAI21X1_202 ( .A(_4917__bF_buf9), .B(_4913__bF_buf4), .C(cpuregs_7_[22]), .Y(_4974_) );
OAI21X1 OAI21X1_203 ( .A(_4824__bF_buf3), .B(_4919__bF_buf2), .C(_4974_), .Y(_144_) );
OAI21X1 OAI21X1_204 ( .A(_4917__bF_buf8), .B(_4913__bF_buf3), .C(cpuregs_7_[23]), .Y(_4975_) );
OAI21X1 OAI21X1_205 ( .A(_4833__bF_buf3), .B(_4919__bF_buf1), .C(_4975_), .Y(_145_) );
OAI21X1 OAI21X1_206 ( .A(_4917__bF_buf7), .B(_4913__bF_buf2), .C(cpuregs_7_[24]), .Y(_4976_) );
OAI21X1 OAI21X1_207 ( .A(_4845__bF_buf3), .B(_4919__bF_buf0), .C(_4976_), .Y(_146_) );
OAI21X1 OAI21X1_208 ( .A(_4917__bF_buf6), .B(_4913__bF_buf1), .C(cpuregs_7_[25]), .Y(_4977_) );
OAI21X1 OAI21X1_209 ( .A(_4854__bF_buf3), .B(_4919__bF_buf4), .C(_4977_), .Y(_147_) );
OAI21X1 OAI21X1_210 ( .A(_4917__bF_buf5), .B(_4913__bF_buf0), .C(cpuregs_7_[26]), .Y(_4978_) );
OAI21X1 OAI21X1_211 ( .A(_4863__bF_buf3), .B(_4919__bF_buf3), .C(_4978_), .Y(_148_) );
OAI21X1 OAI21X1_212 ( .A(_4917__bF_buf4), .B(_4913__bF_buf6), .C(cpuregs_7_[27]), .Y(_4979_) );
OAI21X1 OAI21X1_213 ( .A(_4871__bF_buf3), .B(_4919__bF_buf2), .C(_4979_), .Y(_149_) );
OAI21X1 OAI21X1_214 ( .A(_4917__bF_buf3), .B(_4913__bF_buf5), .C(cpuregs_7_[28]), .Y(_4980_) );
OAI21X1 OAI21X1_215 ( .A(_4884__bF_buf3), .B(_4919__bF_buf1), .C(_4980_), .Y(_150_) );
OAI21X1 OAI21X1_216 ( .A(_4917__bF_buf2), .B(_4913__bF_buf4), .C(cpuregs_7_[29]), .Y(_4981_) );
OAI21X1 OAI21X1_217 ( .A(_4893__bF_buf3), .B(_4919__bF_buf0), .C(_4981_), .Y(_151_) );
OAI21X1 OAI21X1_218 ( .A(_4917__bF_buf1), .B(_4913__bF_buf3), .C(cpuregs_7_[30]), .Y(_4982_) );
OAI21X1 OAI21X1_219 ( .A(_4901__bF_buf3), .B(_4919__bF_buf4), .C(_4982_), .Y(_152_) );
OAI21X1 OAI21X1_220 ( .A(_4917__bF_buf0), .B(_4913__bF_buf2), .C(cpuregs_7_[31]), .Y(_4983_) );
OAI21X1 OAI21X1_221 ( .A(_4910__bF_buf3), .B(_4919__bF_buf3), .C(_4983_), .Y(_153_) );
INVX1 INVX1_156 ( .A(mem_do_rinst_bF_buf0), .Y(_4984_) );
NOR2X1 NOR2X1_122 ( .A(_4984_), .B(_4588_), .Y(_4985_) );
NOR2X1 NOR2X1_123 ( .A(cpu_state_0_), .B(cpu_state_1_bF_buf3_), .Y(_4986_) );
NAND2X1 NAND2X1_80 ( .A(_4445_), .B(_4986_), .Y(_4987_) );
NOR2X1 NOR2X1_124 ( .A(cpu_state_3_bF_buf1_), .B(_4987_), .Y(_4988_) );
AND2X2 AND2X2_13 ( .A(_4589_), .B(_4988_), .Y(_7_) );
NOR2X1 NOR2X1_125 ( .A(_4985__bF_buf8), .B(_7_), .Y(_4989_) );
INVX1 INVX1_157 ( .A(is_slti_blt_slt), .Y(_4990_) );
INVX1 INVX1_158 ( .A(_10734__31_), .Y(_4991_) );
NOR2X1 NOR2X1_126 ( .A(_10735__31_), .B(_4991_), .Y(_4992_) );
NOR2X1 NOR2X1_127 ( .A(_10734__31_), .B(_10735__31_), .Y(_4993_) );
INVX1 INVX1_159 ( .A(_10735__31_), .Y(_4994_) );
NOR2X1 NOR2X1_128 ( .A(_4991_), .B(_4994_), .Y(_4995_) );
NOR2X1 NOR2X1_129 ( .A(_4993_), .B(_4995_), .Y(_4996_) );
INVX1 INVX1_160 ( .A(_4996_), .Y(_4997_) );
INVX1 INVX1_161 ( .A(_10734__30_), .Y(_4998_) );
INVX1 INVX1_162 ( .A(_10735__30_), .Y(_4999_) );
NOR2X1 NOR2X1_130 ( .A(_4998_), .B(_4999_), .Y(_5000_) );
NOR2X1 NOR2X1_131 ( .A(_10734__30_), .B(_10735__30_), .Y(_5001_) );
NOR2X1 NOR2X1_132 ( .A(_5001_), .B(_5000_), .Y(_5002_) );
NOR2X1 NOR2X1_133 ( .A(_4996_), .B(_5002_), .Y(_5003_) );
INVX1 INVX1_163 ( .A(_10734__28_), .Y(_5004_) );
INVX1 INVX1_164 ( .A(_10735__28_), .Y(_5005_) );
NOR2X1 NOR2X1_134 ( .A(_5004_), .B(_5005_), .Y(_5006_) );
NOR2X1 NOR2X1_135 ( .A(_10734__28_), .B(_10735__28_), .Y(_5007_) );
NOR2X1 NOR2X1_136 ( .A(_5007_), .B(_5006_), .Y(_5008_) );
INVX1 INVX1_165 ( .A(_10734__29_), .Y(_5009_) );
INVX1 INVX1_166 ( .A(_10735__29_), .Y(_5010_) );
NOR2X1 NOR2X1_137 ( .A(_5009_), .B(_5010_), .Y(_5011_) );
NOR2X1 NOR2X1_138 ( .A(_10734__29_), .B(_10735__29_), .Y(_5012_) );
NOR2X1 NOR2X1_139 ( .A(_5012_), .B(_5011_), .Y(_5013_) );
NOR2X1 NOR2X1_140 ( .A(_5008_), .B(_5013_), .Y(_5014_) );
NAND2X1 NAND2X1_81 ( .A(_5003_), .B(_5014_), .Y(_5015_) );
INVX1 INVX1_167 ( .A(_10734__27_), .Y(_5016_) );
INVX1 INVX1_168 ( .A(_10735__27_), .Y(_5017_) );
NOR2X1 NOR2X1_141 ( .A(_5016_), .B(_5017_), .Y(_5018_) );
NOR2X1 NOR2X1_142 ( .A(_10734__27_), .B(_10735__27_), .Y(_5019_) );
NOR2X1 NOR2X1_143 ( .A(_5019_), .B(_5018_), .Y(_5020_) );
INVX1 INVX1_169 ( .A(_10734__26_), .Y(_5021_) );
INVX1 INVX1_170 ( .A(_10735__26_), .Y(_5022_) );
NOR2X1 NOR2X1_144 ( .A(_5021_), .B(_5022_), .Y(_5023_) );
NOR2X1 NOR2X1_145 ( .A(_10734__26_), .B(_10735__26_), .Y(_5024_) );
NOR2X1 NOR2X1_146 ( .A(_5024_), .B(_5023_), .Y(_5025_) );
NOR2X1 NOR2X1_147 ( .A(_5020_), .B(_5025_), .Y(_5026_) );
INVX1 INVX1_171 ( .A(_10734__25_), .Y(_5027_) );
INVX1 INVX1_172 ( .A(_10735__25_), .Y(_5028_) );
NOR2X1 NOR2X1_148 ( .A(_5027_), .B(_5028_), .Y(_5029_) );
NOR2X1 NOR2X1_149 ( .A(_10734__25_), .B(_10735__25_), .Y(_5030_) );
NOR2X1 NOR2X1_150 ( .A(_5030_), .B(_5029_), .Y(_5031_) );
INVX1 INVX1_173 ( .A(_10734__24_), .Y(_5032_) );
INVX1 INVX1_174 ( .A(_10735__24_), .Y(_5033_) );
NOR2X1 NOR2X1_151 ( .A(_5032_), .B(_5033_), .Y(_5034_) );
NOR2X1 NOR2X1_152 ( .A(_10734__24_), .B(_10735__24_), .Y(_5035_) );
NOR2X1 NOR2X1_153 ( .A(_5035_), .B(_5034_), .Y(_5036_) );
NOR2X1 NOR2X1_154 ( .A(_5031_), .B(_5036_), .Y(_5037_) );
NAND2X1 NAND2X1_82 ( .A(_5026_), .B(_5037_), .Y(_5038_) );
NOR2X1 NOR2X1_155 ( .A(_5015_), .B(_5038_), .Y(_5039_) );
INVX1 INVX1_175 ( .A(_10734__19_), .Y(_5040_) );
INVX1 INVX1_176 ( .A(_10735__19_), .Y(_5041_) );
NOR2X1 NOR2X1_156 ( .A(_5040_), .B(_5041_), .Y(_5042_) );
NOR2X1 NOR2X1_157 ( .A(_10734__19_), .B(_10735__19_), .Y(_5043_) );
NOR2X1 NOR2X1_158 ( .A(_5043_), .B(_5042_), .Y(_5044_) );
INVX1 INVX1_177 ( .A(_10734__18_), .Y(_5045_) );
INVX1 INVX1_178 ( .A(_10735__18_), .Y(_5046_) );
NOR2X1 NOR2X1_159 ( .A(_5045_), .B(_5046_), .Y(_5047_) );
NOR2X1 NOR2X1_160 ( .A(_10734__18_), .B(_10735__18_), .Y(_5048_) );
NOR2X1 NOR2X1_161 ( .A(_5048_), .B(_5047_), .Y(_5049_) );
NOR2X1 NOR2X1_162 ( .A(_5044_), .B(_5049_), .Y(_5050_) );
INVX1 INVX1_179 ( .A(_10734__16_), .Y(_5051_) );
INVX1 INVX1_180 ( .A(_10735__16_), .Y(_5052_) );
NOR2X1 NOR2X1_163 ( .A(_5051_), .B(_5052_), .Y(_5053_) );
NOR2X1 NOR2X1_164 ( .A(_10734__16_), .B(_10735__16_), .Y(_5054_) );
NOR2X1 NOR2X1_165 ( .A(_5054_), .B(_5053_), .Y(_5055_) );
INVX1 INVX1_181 ( .A(_5055_), .Y(_5056_) );
INVX1 INVX1_182 ( .A(_10734__17_), .Y(_5057_) );
INVX1 INVX1_183 ( .A(_10735__17_), .Y(_5058_) );
NOR2X1 NOR2X1_166 ( .A(_5057_), .B(_5058_), .Y(_5059_) );
NOR2X1 NOR2X1_167 ( .A(_10734__17_), .B(_10735__17_), .Y(_5060_) );
NOR2X1 NOR2X1_168 ( .A(_5060_), .B(_5059_), .Y(_5061_) );
INVX1 INVX1_184 ( .A(_5061_), .Y(_5062_) );
NAND3X1 NAND3X1_17 ( .A(_5056_), .B(_5062_), .C(_5050_), .Y(_5063_) );
NAND2X1 NAND2X1_83 ( .A(_10734__23_), .B(_10735__23_), .Y(_5064_) );
INVX1 INVX1_185 ( .A(_5064_), .Y(_5065_) );
NOR2X1 NOR2X1_169 ( .A(_10734__23_), .B(_10735__23_), .Y(_5066_) );
NOR2X1 NOR2X1_170 ( .A(_5066_), .B(_5065_), .Y(_5067_) );
NAND2X1 NAND2X1_84 ( .A(_10734__22_), .B(_10735__22_), .Y(_5068_) );
INVX1 INVX1_186 ( .A(_5068_), .Y(_5069_) );
NOR2X1 NOR2X1_171 ( .A(_10734__22_), .B(_10735__22_), .Y(_5070_) );
NOR2X1 NOR2X1_172 ( .A(_5070_), .B(_5069_), .Y(_5071_) );
NOR2X1 NOR2X1_173 ( .A(_5067_), .B(_5071_), .Y(_5072_) );
NAND2X1 NAND2X1_85 ( .A(_10734__20_), .B(_10735__20_), .Y(_5073_) );
INVX1 INVX1_187 ( .A(_5073_), .Y(_5074_) );
NOR2X1 NOR2X1_174 ( .A(_10734__20_), .B(_10735__20_), .Y(_5075_) );
NOR2X1 NOR2X1_175 ( .A(_5075_), .B(_5074_), .Y(_5076_) );
NAND2X1 NAND2X1_86 ( .A(_10734__21_), .B(_10735__21_), .Y(_5077_) );
INVX1 INVX1_188 ( .A(_5077_), .Y(_5078_) );
NOR2X1 NOR2X1_176 ( .A(_10734__21_), .B(_10735__21_), .Y(_5079_) );
NOR2X1 NOR2X1_177 ( .A(_5079_), .B(_5078_), .Y(_5080_) );
NOR2X1 NOR2X1_178 ( .A(_5076_), .B(_5080_), .Y(_5081_) );
NAND2X1 NAND2X1_87 ( .A(_5072_), .B(_5081_), .Y(_5082_) );
NOR2X1 NOR2X1_179 ( .A(_5082_), .B(_5063_), .Y(_5083_) );
NAND2X1 NAND2X1_88 ( .A(_5039_), .B(_5083_), .Y(_5084_) );
INVX1 INVX1_189 ( .A(_5084_), .Y(_5085_) );
NAND2X1 NAND2X1_89 ( .A(_10734__15_), .B(_10735__15_), .Y(_5086_) );
INVX1 INVX1_190 ( .A(_10734__15_), .Y(_5087_) );
INVX1 INVX1_191 ( .A(_10735__15_), .Y(_5088_) );
NAND2X1 NAND2X1_90 ( .A(_5087_), .B(_5088_), .Y(_5089_) );
NAND2X1 NAND2X1_91 ( .A(_5086_), .B(_5089_), .Y(_5090_) );
NAND2X1 NAND2X1_92 ( .A(_10734__14_), .B(_10735__14_), .Y(_5091_) );
INVX1 INVX1_192 ( .A(_5091_), .Y(_5092_) );
NOR2X1 NOR2X1_180 ( .A(_10734__14_), .B(_10735__14_), .Y(_5093_) );
OAI21X1 OAI21X1_222 ( .A(_5092_), .B(_5093_), .C(_5090_), .Y(_5094_) );
NAND2X1 NAND2X1_93 ( .A(_10734__12_), .B(_10735__12_), .Y(_5095_) );
INVX1 INVX1_193 ( .A(_5095_), .Y(_5096_) );
NOR2X1 NOR2X1_181 ( .A(_10734__12_), .B(_10735__12_), .Y(_5097_) );
NOR2X1 NOR2X1_182 ( .A(_5097_), .B(_5096_), .Y(_5098_) );
INVX1 INVX1_194 ( .A(_5098_), .Y(_5099_) );
NAND2X1 NAND2X1_94 ( .A(_10734__13_), .B(_10735__13_), .Y(_5100_) );
INVX1 INVX1_195 ( .A(_5100_), .Y(_5101_) );
NOR2X1 NOR2X1_183 ( .A(_10734__13_), .B(_10735__13_), .Y(_5102_) );
OAI21X1 OAI21X1_223 ( .A(_5101_), .B(_5102_), .C(_5099_), .Y(_5103_) );
NOR2X1 NOR2X1_184 ( .A(_5094_), .B(_5103_), .Y(_5104_) );
INVX1 INVX1_196 ( .A(_5104_), .Y(_5105_) );
NOR2X1 NOR2X1_185 ( .A(_10734__9_), .B(_10735__9_), .Y(_5106_) );
INVX1 INVX1_197 ( .A(_10734__9_), .Y(_5107_) );
INVX1 INVX1_198 ( .A(_10735__9_), .Y(_5108_) );
NOR2X1 NOR2X1_186 ( .A(_5107_), .B(_5108_), .Y(_5109_) );
NAND2X1 NAND2X1_95 ( .A(_10734__8_), .B(_10735__8_), .Y(_5110_) );
INVX1 INVX1_199 ( .A(_5110_), .Y(_5111_) );
NOR2X1 NOR2X1_187 ( .A(_10734__8_), .B(_10735__8_), .Y(_5112_) );
NOR2X1 NOR2X1_188 ( .A(_5112_), .B(_5111_), .Y(_5113_) );
INVX1 INVX1_200 ( .A(_5113_), .Y(_5114_) );
OAI21X1 OAI21X1_224 ( .A(_5106_), .B(_5109_), .C(_5114_), .Y(_5115_) );
NAND2X1 NAND2X1_96 ( .A(_10734__11_), .B(_10735__11_), .Y(_5116_) );
INVX1 INVX1_201 ( .A(_10734__11_), .Y(_5117_) );
INVX1 INVX1_202 ( .A(_10735__11_), .Y(_5118_) );
NAND2X1 NAND2X1_97 ( .A(_5117_), .B(_5118_), .Y(_5119_) );
NAND2X1 NAND2X1_98 ( .A(_5116_), .B(_5119_), .Y(_5120_) );
INVX1 INVX1_203 ( .A(_10734__10_), .Y(_5121_) );
INVX1 INVX1_204 ( .A(_10735__10_), .Y(_5122_) );
NOR2X1 NOR2X1_189 ( .A(_5121_), .B(_5122_), .Y(_5123_) );
NOR2X1 NOR2X1_190 ( .A(_10734__10_), .B(_10735__10_), .Y(_5124_) );
OAI21X1 OAI21X1_225 ( .A(_5123_), .B(_5124_), .C(_5120_), .Y(_5125_) );
NOR2X1 NOR2X1_191 ( .A(_5125_), .B(_5115_), .Y(_5126_) );
INVX1 INVX1_205 ( .A(_5126_), .Y(_5127_) );
NOR2X1 NOR2X1_192 ( .A(_5105_), .B(_5127_), .Y(_5128_) );
INVX1 INVX1_206 ( .A(_5128_), .Y(_5129_) );
INVX1 INVX1_207 ( .A(_10734__3_), .Y(_5130_) );
INVX1 INVX1_208 ( .A(_10728__2_bF_buf4_), .Y(_5131_) );
NAND2X1 NAND2X1_99 ( .A(_10734__2_), .B(_5131__bF_buf5), .Y(_5132_) );
NAND2X1 NAND2X1_100 ( .A(_10734__3_), .B(_10728__3_bF_buf4_), .Y(_5133_) );
NOR2X1 NOR2X1_193 ( .A(_10734__3_), .B(_10728__3_bF_buf3_), .Y(_5134_) );
INVX1 INVX1_209 ( .A(_5134_), .Y(_5135_) );
NAND2X1 NAND2X1_101 ( .A(_5133_), .B(_5135_), .Y(_5136_) );
INVX1 INVX1_210 ( .A(_5136_), .Y(_5137_) );
OR2X2 OR2X2_2 ( .A(_5137_), .B(_5132_), .Y(_5138_) );
OAI21X1 OAI21X1_226 ( .A(_5130_), .B(_10728__3_bF_buf2_), .C(_5138_), .Y(_5139_) );
INVX1 INVX1_211 ( .A(_10728__1_bF_buf3_), .Y(_5140_) );
NAND2X1 NAND2X1_102 ( .A(_10734__1_), .B(_5140__bF_buf5), .Y(_5141_) );
INVX1 INVX1_212 ( .A(_10728__0_bF_buf7_), .Y(_5142_) );
NAND2X1 NAND2X1_103 ( .A(_10734__1_), .B(_10728__1_bF_buf2_), .Y(_5143_) );
NAND2X1 NAND2X1_104 ( .A(_4490_), .B(_5140__bF_buf4), .Y(_5144_) );
NAND2X1 NAND2X1_105 ( .A(_5143_), .B(_5144_), .Y(_5145_) );
OAI21X1 OAI21X1_227 ( .A(_10734__0_), .B(_5142_), .C(_5145_), .Y(_5146_) );
AND2X2 AND2X2_14 ( .A(_5146_), .B(_5141_), .Y(_5147_) );
INVX1 INVX1_213 ( .A(_10734__2_), .Y(_5148_) );
NOR2X1 NOR2X1_194 ( .A(_5148_), .B(_5131__bF_buf4), .Y(_5149_) );
NOR2X1 NOR2X1_195 ( .A(_10734__2_), .B(_10728__2_bF_buf3_), .Y(_5150_) );
OAI21X1 OAI21X1_228 ( .A(_5149_), .B(_5150_), .C(_5136_), .Y(_5151_) );
NOR2X1 NOR2X1_196 ( .A(_5151_), .B(_5147_), .Y(_5152_) );
NAND2X1 NAND2X1_106 ( .A(_10734__7_), .B(_10728__7_), .Y(_5153_) );
INVX1 INVX1_214 ( .A(_5153_), .Y(_5154_) );
NOR2X1 NOR2X1_197 ( .A(_10734__7_), .B(_10728__7_), .Y(_5155_) );
NOR2X1 NOR2X1_198 ( .A(_5155_), .B(_5154_), .Y(_5156_) );
INVX1 INVX1_215 ( .A(_5156_), .Y(_5157_) );
NAND2X1 NAND2X1_107 ( .A(_10734__6_), .B(_10728__6_), .Y(_5158_) );
INVX1 INVX1_216 ( .A(_5158_), .Y(_5159_) );
NOR2X1 NOR2X1_199 ( .A(_10734__6_), .B(_10728__6_), .Y(_5160_) );
OAI21X1 OAI21X1_229 ( .A(_5159_), .B(_5160_), .C(_5157_), .Y(_5161_) );
NOR2X1 NOR2X1_200 ( .A(_10734__5_), .B(_10728__5_), .Y(_5162_) );
NAND2X1 NAND2X1_108 ( .A(_10734__5_), .B(_10728__5_), .Y(_5163_) );
INVX1 INVX1_217 ( .A(_5163_), .Y(_5164_) );
NOR2X1 NOR2X1_201 ( .A(_5162_), .B(_5164_), .Y(_5165_) );
INVX1 INVX1_218 ( .A(_5165_), .Y(_5166_) );
NAND2X1 NAND2X1_109 ( .A(_10734__4_), .B(_10728__4_bF_buf4_), .Y(_5167_) );
INVX1 INVX1_219 ( .A(_5167_), .Y(_5168_) );
NOR2X1 NOR2X1_202 ( .A(_10734__4_), .B(_10728__4_bF_buf3_), .Y(_5169_) );
OAI21X1 OAI21X1_230 ( .A(_5168_), .B(_5169_), .C(_5166_), .Y(_5170_) );
NOR2X1 NOR2X1_203 ( .A(_5161_), .B(_5170_), .Y(_5171_) );
OAI21X1 OAI21X1_231 ( .A(_5152_), .B(_5139_), .C(_5171_), .Y(_5172_) );
INVX1 INVX1_220 ( .A(_10734__7_), .Y(_5173_) );
INVX1 INVX1_221 ( .A(_10734__6_), .Y(_5174_) );
NOR2X1 NOR2X1_204 ( .A(_10728__6_), .B(_5174_), .Y(_5175_) );
OAI21X1 OAI21X1_232 ( .A(_5154_), .B(_5155_), .C(_5175_), .Y(_5176_) );
OAI21X1 OAI21X1_233 ( .A(_5173_), .B(_10728__7_), .C(_5176_), .Y(_5177_) );
INVX1 INVX1_222 ( .A(_5161_), .Y(_5178_) );
INVX1 INVX1_223 ( .A(_10734__5_), .Y(_5179_) );
INVX1 INVX1_224 ( .A(_10734__4_), .Y(_5180_) );
NOR2X1 NOR2X1_205 ( .A(_10728__4_bF_buf2_), .B(_5180_), .Y(_5181_) );
OAI21X1 OAI21X1_234 ( .A(_5164_), .B(_5162_), .C(_5181_), .Y(_5182_) );
OAI21X1 OAI21X1_235 ( .A(_5179_), .B(_10728__5_), .C(_5182_), .Y(_5183_) );
AOI21X1 AOI21X1_13 ( .A(_5183_), .B(_5178_), .C(_5177_), .Y(_5184_) );
AND2X2 AND2X2_15 ( .A(_5172_), .B(_5184_), .Y(_5185_) );
NOR2X1 NOR2X1_206 ( .A(_5129_), .B(_5185_), .Y(_5186_) );
INVX1 INVX1_225 ( .A(_10734__8_), .Y(_5187_) );
NOR2X1 NOR2X1_207 ( .A(_10735__8_), .B(_5187_), .Y(_5188_) );
OAI21X1 OAI21X1_236 ( .A(_5109_), .B(_5106_), .C(_5188_), .Y(_5189_) );
NAND2X1 NAND2X1_110 ( .A(_10734__9_), .B(_5108_), .Y(_5190_) );
AND2X2 AND2X2_16 ( .A(_5189_), .B(_5190_), .Y(_5191_) );
NAND3X1 NAND3X1_18 ( .A(_10734__10_), .B(_5122_), .C(_5120_), .Y(_5192_) );
OAI21X1 OAI21X1_237 ( .A(_5191_), .B(_5125_), .C(_5192_), .Y(_5193_) );
AOI21X1 AOI21X1_14 ( .A(_10734__11_), .B(_5118_), .C(_5193_), .Y(_5194_) );
NOR2X1 NOR2X1_208 ( .A(_5105_), .B(_5194_), .Y(_5195_) );
INVX1 INVX1_226 ( .A(_10734__13_), .Y(_5196_) );
INVX1 INVX1_227 ( .A(_10734__12_), .Y(_5197_) );
NOR2X1 NOR2X1_209 ( .A(_10735__12_), .B(_5197_), .Y(_5198_) );
OAI21X1 OAI21X1_238 ( .A(_5101_), .B(_5102_), .C(_5198_), .Y(_5199_) );
OAI21X1 OAI21X1_239 ( .A(_5196_), .B(_10735__13_), .C(_5199_), .Y(_5200_) );
INVX1 INVX1_228 ( .A(_5200_), .Y(_5201_) );
NOR2X1 NOR2X1_210 ( .A(_10735__15_), .B(_5087_), .Y(_5202_) );
INVX1 INVX1_229 ( .A(_10734__14_), .Y(_5203_) );
NOR2X1 NOR2X1_211 ( .A(_10735__14_), .B(_5203_), .Y(_5204_) );
AOI21X1 AOI21X1_15 ( .A(_5204_), .B(_5090_), .C(_5202_), .Y(_5205_) );
OAI21X1 OAI21X1_240 ( .A(_5201_), .B(_5094_), .C(_5205_), .Y(_5206_) );
OR2X2 OR2X2_3 ( .A(_5195_), .B(_5206_), .Y(_5207_) );
OAI21X1 OAI21X1_241 ( .A(_5186_), .B(_5207_), .C(_5085_), .Y(_5208_) );
NAND2X1 NAND2X1_111 ( .A(_10734__16_), .B(_5052_), .Y(_5209_) );
NAND2X1 NAND2X1_112 ( .A(_10734__17_), .B(_5058_), .Y(_5210_) );
OAI21X1 OAI21X1_242 ( .A(_5061_), .B(_5209_), .C(_5210_), .Y(_5211_) );
INVX1 INVX1_230 ( .A(_5044_), .Y(_5212_) );
NAND3X1 NAND3X1_19 ( .A(_10734__18_), .B(_5046_), .C(_5212_), .Y(_5213_) );
OAI21X1 OAI21X1_243 ( .A(_5040_), .B(_10735__19_), .C(_5213_), .Y(_5214_) );
AOI21X1 AOI21X1_16 ( .A(_5050_), .B(_5211_), .C(_5214_), .Y(_5215_) );
NOR2X1 NOR2X1_212 ( .A(_5082_), .B(_5215_), .Y(_5216_) );
INVX1 INVX1_231 ( .A(_10734__21_), .Y(_5217_) );
INVX1 INVX1_232 ( .A(_10734__20_), .Y(_5218_) );
NOR2X1 NOR2X1_213 ( .A(_10735__20_), .B(_5218_), .Y(_5219_) );
OAI21X1 OAI21X1_244 ( .A(_5078_), .B(_5079_), .C(_5219_), .Y(_5220_) );
OAI21X1 OAI21X1_245 ( .A(_5217_), .B(_10735__21_), .C(_5220_), .Y(_5221_) );
NAND2X1 NAND2X1_113 ( .A(_5221_), .B(_5072_), .Y(_5222_) );
INVX1 INVX1_233 ( .A(_10735__23_), .Y(_5223_) );
INVX1 INVX1_234 ( .A(_10735__22_), .Y(_5224_) );
NAND2X1 NAND2X1_114 ( .A(_10734__22_), .B(_5224_), .Y(_5225_) );
NOR2X1 NOR2X1_214 ( .A(_5225_), .B(_5067_), .Y(_5226_) );
AOI21X1 AOI21X1_17 ( .A(_10734__23_), .B(_5223_), .C(_5226_), .Y(_5227_) );
NAND2X1 NAND2X1_115 ( .A(_5222_), .B(_5227_), .Y(_5228_) );
OR2X2 OR2X2_4 ( .A(_5216_), .B(_5228_), .Y(_5229_) );
NOR2X1 NOR2X1_215 ( .A(_10735__24_), .B(_5032_), .Y(_5230_) );
OAI21X1 OAI21X1_246 ( .A(_5029_), .B(_5030_), .C(_5230_), .Y(_5231_) );
OAI21X1 OAI21X1_247 ( .A(_5027_), .B(_10735__25_), .C(_5231_), .Y(_5232_) );
NAND2X1 NAND2X1_116 ( .A(_5232_), .B(_5026_), .Y(_5233_) );
INVX1 INVX1_235 ( .A(_5233_), .Y(_5234_) );
NOR2X1 NOR2X1_216 ( .A(_10735__26_), .B(_5021_), .Y(_5235_) );
OAI21X1 OAI21X1_248 ( .A(_5018_), .B(_5019_), .C(_5235_), .Y(_5236_) );
OAI21X1 OAI21X1_249 ( .A(_5016_), .B(_10735__27_), .C(_5236_), .Y(_5237_) );
OR2X2 OR2X2_5 ( .A(_5234_), .B(_5237_), .Y(_5238_) );
INVX1 INVX1_236 ( .A(_5238_), .Y(_5239_) );
NOR2X1 NOR2X1_217 ( .A(_10735__28_), .B(_5004_), .Y(_5240_) );
OAI21X1 OAI21X1_250 ( .A(_5011_), .B(_5012_), .C(_5240_), .Y(_5241_) );
OAI21X1 OAI21X1_251 ( .A(_5009_), .B(_10735__29_), .C(_5241_), .Y(_5242_) );
NOR2X1 NOR2X1_218 ( .A(_10735__30_), .B(_4998_), .Y(_5243_) );
OAI21X1 OAI21X1_252 ( .A(_4995_), .B(_4993_), .C(_5243_), .Y(_5244_) );
OAI21X1 OAI21X1_253 ( .A(_4991_), .B(_10735__31_), .C(_5244_), .Y(_5245_) );
AOI21X1 AOI21X1_18 ( .A(_5242_), .B(_5003_), .C(_5245_), .Y(_5246_) );
OAI21X1 OAI21X1_254 ( .A(_5239_), .B(_5015_), .C(_5246_), .Y(_5247_) );
AOI21X1 AOI21X1_19 ( .A(_5039_), .B(_5229_), .C(_5247_), .Y(_5248_) );
AND2X2 AND2X2_17 ( .A(_5208_), .B(_5248_), .Y(_5249_) );
AOI21X1 AOI21X1_20 ( .A(_4997_), .B(_5249_), .C(_4992_), .Y(_5250_) );
NOR2X1 NOR2X1_219 ( .A(_4990_), .B(_5250_), .Y(_5251_) );
INVX1 INVX1_237 ( .A(instr_bgeu), .Y(_5252_) );
NAND2X1 NAND2X1_117 ( .A(_10734__0_), .B(_10728__0_bF_buf6_), .Y(_5253_) );
INVX1 INVX1_238 ( .A(_5253_), .Y(_5254_) );
NOR2X1 NOR2X1_220 ( .A(_10734__0_), .B(_10728__0_bF_buf5_), .Y(_5255_) );
OAI21X1 OAI21X1_255 ( .A(_5254_), .B(_5255_), .C(_5145_), .Y(_5256_) );
NOR2X1 NOR2X1_221 ( .A(_5256_), .B(_5151_), .Y(_5257_) );
NAND3X1 NAND3X1_20 ( .A(_5171_), .B(_5257_), .C(_5128_), .Y(_5258_) );
NOR2X1 NOR2X1_222 ( .A(_5084_), .B(_5258_), .Y(_5259_) );
MUX2X1 MUX2X1_14 ( .A(instr_beq), .B(instr_bne), .S(_5259_), .Y(_5260_) );
OAI21X1 OAI21X1_256 ( .A(_5249_), .B(_5252_), .C(_5260_), .Y(_5261_) );
NAND2X1 NAND2X1_118 ( .A(instr_bge), .B(_5250_), .Y(_5262_) );
NOR2X1 NOR2X1_223 ( .A(is_slti_blt_slt), .B(_4507_), .Y(_5263_) );
NAND2X1 NAND2X1_119 ( .A(_5263_), .B(_5249_), .Y(_5264_) );
NAND2X1 NAND2X1_120 ( .A(_5264_), .B(_5262_), .Y(_5265_) );
NOR3X1 NOR3X1_1 ( .A(_5251_), .B(_5261_), .C(_5265_), .Y(_5266_) );
OAI21X1 OAI21X1_257 ( .A(_5266_), .B(_4556_), .C(cpu_state_3_bF_buf0_), .Y(_5267_) );
NOR2X1 NOR2X1_224 ( .A(_4555_), .B(_4987_), .Y(_5268_) );
AOI21X1 AOI21X1_21 ( .A(_5268_), .B(_5267_), .C(_4989_), .Y(_8_) );
INVX1 INVX1_239 ( .A(cpuregs_6_[0]), .Y(_5269_) );
NOR2X1 NOR2X1_225 ( .A(latched_rd_0_), .B(_4914_), .Y(_5270_) );
NAND2X1 NAND2X1_121 ( .A(_5270_), .B(_4912_), .Y(_5271_) );
NOR2X1 NOR2X1_226 ( .A(_5271__bF_buf3), .B(_4632__bF_buf5), .Y(_5272_) );
INVX1 INVX1_240 ( .A(_4925__bF_buf3), .Y(_5273_) );
NAND2X1 NAND2X1_122 ( .A(_5273_), .B(_5272_), .Y(_5274_) );
OAI21X1 OAI21X1_258 ( .A(_5269_), .B(_5272_), .C(_5274_), .Y(_154_) );
INVX1 INVX1_241 ( .A(cpuregs_6_[1]), .Y(_5275_) );
MUX2X1 MUX2X1_15 ( .A(_4933__bF_buf3), .B(_5275_), .S(_5272_), .Y(_155_) );
INVX1 INVX1_242 ( .A(cpuregs_6_[2]), .Y(_5276_) );
MUX2X1 MUX2X1_16 ( .A(_4940__bF_buf3), .B(_5276_), .S(_5272_), .Y(_156_) );
INVX1 INVX1_243 ( .A(cpuregs_6_[3]), .Y(_5277_) );
MUX2X1 MUX2X1_17 ( .A(_4948__bF_buf3), .B(_5277_), .S(_5272_), .Y(_157_) );
INVX1 INVX1_244 ( .A(cpuregs_6_[4]), .Y(_5278_) );
INVX1 INVX1_245 ( .A(_4955__bF_buf3), .Y(_5279_) );
NAND2X1 NAND2X1_123 ( .A(_5272_), .B(_5279_), .Y(_5280_) );
OAI21X1 OAI21X1_259 ( .A(_5278_), .B(_5272_), .C(_5280_), .Y(_158_) );
NAND2X1 NAND2X1_124 ( .A(_5270_), .B(_4631_), .Y(_5281_) );
NOR2X1 NOR2X1_227 ( .A(_4913__bF_buf1), .B(_5281__bF_buf10), .Y(_5282_) );
NOR2X1 NOR2X1_228 ( .A(cpuregs_6_[5]), .B(_5282_), .Y(_5283_) );
AOI21X1 AOI21X1_22 ( .A(_4654__bF_buf2), .B(_5282_), .C(_5283_), .Y(_159_) );
NOR2X1 NOR2X1_229 ( .A(cpuregs_6_[6]), .B(_5282_), .Y(_5284_) );
AOI21X1 AOI21X1_23 ( .A(_5282_), .B(_4664__bF_buf2), .C(_5284_), .Y(_160_) );
NOR2X1 NOR2X1_230 ( .A(cpuregs_6_[7]), .B(_5282_), .Y(_5285_) );
AOI21X1 AOI21X1_24 ( .A(_5282_), .B(_4677__bF_buf2), .C(_5285_), .Y(_161_) );
NOR2X1 NOR2X1_231 ( .A(cpuregs_6_[8]), .B(_5282_), .Y(_5286_) );
AOI21X1 AOI21X1_25 ( .A(_5282_), .B(_4685__bF_buf2), .C(_5286_), .Y(_162_) );
NOR2X1 NOR2X1_232 ( .A(cpuregs_6_[9]), .B(_5282_), .Y(_5287_) );
AOI21X1 AOI21X1_26 ( .A(_5282_), .B(_4696__bF_buf2), .C(_5287_), .Y(_163_) );
NOR2X1 NOR2X1_233 ( .A(cpuregs_6_[10]), .B(_5282_), .Y(_5288_) );
AOI21X1 AOI21X1_27 ( .A(_5282_), .B(_4703__bF_buf2), .C(_5288_), .Y(_164_) );
INVX1 INVX1_246 ( .A(cpuregs_6_[11]), .Y(_5289_) );
MUX2X1 MUX2X1_18 ( .A(_4713__bF_buf2), .B(_5289_), .S(_5282_), .Y(_165_) );
INVX1 INVX1_247 ( .A(_5282_), .Y(_5290_) );
OAI21X1 OAI21X1_260 ( .A(_4632__bF_buf4), .B(_5271__bF_buf2), .C(cpuregs_6_[12]), .Y(_5291_) );
OAI21X1 OAI21X1_261 ( .A(_4722__bF_buf2), .B(_5290__bF_buf3), .C(_5291_), .Y(_166_) );
OAI21X1 OAI21X1_262 ( .A(_4632__bF_buf3), .B(_5271__bF_buf1), .C(cpuregs_6_[13]), .Y(_5292_) );
OAI21X1 OAI21X1_263 ( .A(_4731__bF_buf2), .B(_5290__bF_buf2), .C(_5292_), .Y(_167_) );
OAI21X1 OAI21X1_264 ( .A(_4632__bF_buf2), .B(_5271__bF_buf0), .C(cpuregs_6_[14]), .Y(_5293_) );
OAI21X1 OAI21X1_265 ( .A(_4740__bF_buf2), .B(_5290__bF_buf1), .C(_5293_), .Y(_168_) );
OAI21X1 OAI21X1_266 ( .A(_4632__bF_buf1), .B(_5271__bF_buf3), .C(cpuregs_6_[15]), .Y(_5294_) );
OAI21X1 OAI21X1_267 ( .A(_4747__bF_buf2), .B(_5290__bF_buf0), .C(_5294_), .Y(_169_) );
OAI21X1 OAI21X1_268 ( .A(_4632__bF_buf0), .B(_5271__bF_buf2), .C(cpuregs_6_[16]), .Y(_5295_) );
OAI21X1 OAI21X1_269 ( .A(_4755__bF_buf2), .B(_5290__bF_buf3), .C(_5295_), .Y(_170_) );
OAI21X1 OAI21X1_270 ( .A(_4632__bF_buf8), .B(_5271__bF_buf1), .C(cpuregs_6_[17]), .Y(_5296_) );
OAI21X1 OAI21X1_271 ( .A(_4763__bF_buf2), .B(_5290__bF_buf2), .C(_5296_), .Y(_171_) );
OAI21X1 OAI21X1_272 ( .A(_4632__bF_buf7), .B(_5271__bF_buf0), .C(cpuregs_6_[18]), .Y(_5297_) );
OAI21X1 OAI21X1_273 ( .A(_4783__bF_buf2), .B(_5290__bF_buf1), .C(_5297_), .Y(_172_) );
OAI21X1 OAI21X1_274 ( .A(_4632__bF_buf6), .B(_5271__bF_buf3), .C(cpuregs_6_[19]), .Y(_5298_) );
OAI21X1 OAI21X1_275 ( .A(_4793__bF_buf2), .B(_5290__bF_buf0), .C(_5298_), .Y(_173_) );
OAI21X1 OAI21X1_276 ( .A(_4632__bF_buf5), .B(_5271__bF_buf2), .C(cpuregs_6_[20]), .Y(_5299_) );
OAI21X1 OAI21X1_277 ( .A(_4806__bF_buf2), .B(_5290__bF_buf3), .C(_5299_), .Y(_174_) );
OAI21X1 OAI21X1_278 ( .A(_4632__bF_buf4), .B(_5271__bF_buf1), .C(cpuregs_6_[21]), .Y(_5300_) );
OAI21X1 OAI21X1_279 ( .A(_4816__bF_buf2), .B(_5290__bF_buf2), .C(_5300_), .Y(_175_) );
OAI21X1 OAI21X1_280 ( .A(_4632__bF_buf3), .B(_5271__bF_buf0), .C(cpuregs_6_[22]), .Y(_5301_) );
OAI21X1 OAI21X1_281 ( .A(_4824__bF_buf2), .B(_5290__bF_buf1), .C(_5301_), .Y(_176_) );
OAI21X1 OAI21X1_282 ( .A(_4632__bF_buf2), .B(_5271__bF_buf3), .C(cpuregs_6_[23]), .Y(_5302_) );
OAI21X1 OAI21X1_283 ( .A(_4833__bF_buf2), .B(_5290__bF_buf0), .C(_5302_), .Y(_177_) );
OAI21X1 OAI21X1_284 ( .A(_4632__bF_buf1), .B(_5271__bF_buf2), .C(cpuregs_6_[24]), .Y(_5303_) );
OAI21X1 OAI21X1_285 ( .A(_4845__bF_buf2), .B(_5290__bF_buf3), .C(_5303_), .Y(_178_) );
OAI21X1 OAI21X1_286 ( .A(_4632__bF_buf0), .B(_5271__bF_buf1), .C(cpuregs_6_[25]), .Y(_5304_) );
OAI21X1 OAI21X1_287 ( .A(_4854__bF_buf2), .B(_5290__bF_buf2), .C(_5304_), .Y(_179_) );
OAI21X1 OAI21X1_288 ( .A(_4632__bF_buf8), .B(_5271__bF_buf0), .C(cpuregs_6_[26]), .Y(_5305_) );
OAI21X1 OAI21X1_289 ( .A(_4863__bF_buf2), .B(_5290__bF_buf1), .C(_5305_), .Y(_180_) );
OAI21X1 OAI21X1_290 ( .A(_4632__bF_buf7), .B(_5271__bF_buf3), .C(cpuregs_6_[27]), .Y(_5306_) );
OAI21X1 OAI21X1_291 ( .A(_4871__bF_buf2), .B(_5290__bF_buf0), .C(_5306_), .Y(_181_) );
OAI21X1 OAI21X1_292 ( .A(_4632__bF_buf6), .B(_5271__bF_buf2), .C(cpuregs_6_[28]), .Y(_5307_) );
OAI21X1 OAI21X1_293 ( .A(_4884__bF_buf2), .B(_5290__bF_buf3), .C(_5307_), .Y(_182_) );
OAI21X1 OAI21X1_294 ( .A(_4632__bF_buf5), .B(_5271__bF_buf1), .C(cpuregs_6_[29]), .Y(_5308_) );
OAI21X1 OAI21X1_295 ( .A(_4893__bF_buf2), .B(_5290__bF_buf2), .C(_5308_), .Y(_183_) );
OAI21X1 OAI21X1_296 ( .A(_4632__bF_buf4), .B(_5271__bF_buf0), .C(cpuregs_6_[30]), .Y(_5309_) );
OAI21X1 OAI21X1_297 ( .A(_4901__bF_buf2), .B(_5290__bF_buf1), .C(_5309_), .Y(_184_) );
OAI21X1 OAI21X1_298 ( .A(_4632__bF_buf3), .B(_5271__bF_buf3), .C(cpuregs_6_[31]), .Y(_5310_) );
OAI21X1 OAI21X1_299 ( .A(_4910__bF_buf2), .B(_5290__bF_buf0), .C(_5310_), .Y(_185_) );
NOR2X1 NOR2X1_234 ( .A(latched_rd_1_), .B(_4915_), .Y(_5311_) );
INVX1 INVX1_248 ( .A(_5311_), .Y(_5312_) );
NOR2X1 NOR2X1_235 ( .A(_5312_), .B(_4632__bF_buf2), .Y(_5313_) );
NAND2X1 NAND2X1_125 ( .A(_4912_), .B(_5313_), .Y(_5314_) );
NAND2X1 NAND2X1_126 ( .A(cpuregs_5_[0]), .B(_5314__bF_buf7), .Y(_5315_) );
OAI21X1 OAI21X1_300 ( .A(_4925__bF_buf2), .B(_5314__bF_buf6), .C(_5315_), .Y(_186_) );
NAND2X1 NAND2X1_127 ( .A(cpuregs_5_[1]), .B(_5314__bF_buf5), .Y(_5316_) );
OAI21X1 OAI21X1_301 ( .A(_4933__bF_buf2), .B(_5314__bF_buf4), .C(_5316_), .Y(_187_) );
NAND2X1 NAND2X1_128 ( .A(cpuregs_5_[2]), .B(_5314__bF_buf3), .Y(_5317_) );
OAI21X1 OAI21X1_302 ( .A(_4940__bF_buf2), .B(_5314__bF_buf2), .C(_5317_), .Y(_188_) );
NAND2X1 NAND2X1_129 ( .A(cpuregs_5_[3]), .B(_5314__bF_buf1), .Y(_5318_) );
OAI21X1 OAI21X1_303 ( .A(_4948__bF_buf2), .B(_5314__bF_buf0), .C(_5318_), .Y(_189_) );
NAND2X1 NAND2X1_130 ( .A(cpuregs_5_[4]), .B(_5314__bF_buf7), .Y(_5319_) );
OAI21X1 OAI21X1_304 ( .A(_4955__bF_buf2), .B(_5314__bF_buf6), .C(_5319_), .Y(_190_) );
NAND2X1 NAND2X1_131 ( .A(cpuregs_5_[5]), .B(_5314__bF_buf5), .Y(_5320_) );
OAI21X1 OAI21X1_305 ( .A(_4654__bF_buf1), .B(_5314__bF_buf4), .C(_5320_), .Y(_191_) );
NAND2X1 NAND2X1_132 ( .A(cpuregs_5_[6]), .B(_5314__bF_buf3), .Y(_5321_) );
OAI21X1 OAI21X1_306 ( .A(_4664__bF_buf1), .B(_5314__bF_buf2), .C(_5321_), .Y(_192_) );
NAND2X1 NAND2X1_133 ( .A(cpuregs_5_[7]), .B(_5314__bF_buf1), .Y(_5322_) );
OAI21X1 OAI21X1_307 ( .A(_4677__bF_buf1), .B(_5314__bF_buf0), .C(_5322_), .Y(_193_) );
NAND2X1 NAND2X1_134 ( .A(cpuregs_5_[8]), .B(_5314__bF_buf7), .Y(_5323_) );
OAI21X1 OAI21X1_308 ( .A(_4685__bF_buf1), .B(_5314__bF_buf6), .C(_5323_), .Y(_194_) );
NAND2X1 NAND2X1_135 ( .A(cpuregs_5_[9]), .B(_5314__bF_buf5), .Y(_5324_) );
OAI21X1 OAI21X1_309 ( .A(_4696__bF_buf1), .B(_5314__bF_buf4), .C(_5324_), .Y(_195_) );
NAND2X1 NAND2X1_136 ( .A(cpuregs_5_[10]), .B(_5314__bF_buf3), .Y(_5325_) );
OAI21X1 OAI21X1_310 ( .A(_4703__bF_buf1), .B(_5314__bF_buf2), .C(_5325_), .Y(_196_) );
NAND2X1 NAND2X1_137 ( .A(cpuregs_5_[11]), .B(_5314__bF_buf1), .Y(_5326_) );
OAI21X1 OAI21X1_311 ( .A(_4713__bF_buf1), .B(_5314__bF_buf0), .C(_5326_), .Y(_197_) );
NAND2X1 NAND2X1_138 ( .A(cpuregs_5_[12]), .B(_5314__bF_buf7), .Y(_5327_) );
OAI21X1 OAI21X1_312 ( .A(_4722__bF_buf1), .B(_5314__bF_buf6), .C(_5327_), .Y(_198_) );
NAND2X1 NAND2X1_139 ( .A(cpuregs_5_[13]), .B(_5314__bF_buf5), .Y(_5328_) );
OAI21X1 OAI21X1_313 ( .A(_4731__bF_buf1), .B(_5314__bF_buf4), .C(_5328_), .Y(_199_) );
NAND2X1 NAND2X1_140 ( .A(cpuregs_5_[14]), .B(_5314__bF_buf3), .Y(_5329_) );
OAI21X1 OAI21X1_314 ( .A(_4740__bF_buf1), .B(_5314__bF_buf2), .C(_5329_), .Y(_200_) );
NAND2X1 NAND2X1_141 ( .A(cpuregs_5_[15]), .B(_5314__bF_buf1), .Y(_5330_) );
OAI21X1 OAI21X1_315 ( .A(_4747__bF_buf1), .B(_5314__bF_buf0), .C(_5330_), .Y(_201_) );
NAND2X1 NAND2X1_142 ( .A(cpuregs_5_[16]), .B(_5314__bF_buf7), .Y(_5331_) );
OAI21X1 OAI21X1_316 ( .A(_4755__bF_buf1), .B(_5314__bF_buf6), .C(_5331_), .Y(_202_) );
NAND2X1 NAND2X1_143 ( .A(cpuregs_5_[17]), .B(_5314__bF_buf5), .Y(_5332_) );
OAI21X1 OAI21X1_317 ( .A(_4763__bF_buf1), .B(_5314__bF_buf4), .C(_5332_), .Y(_203_) );
NAND2X1 NAND2X1_144 ( .A(cpuregs_5_[18]), .B(_5314__bF_buf3), .Y(_5333_) );
OAI21X1 OAI21X1_318 ( .A(_4783__bF_buf1), .B(_5314__bF_buf2), .C(_5333_), .Y(_204_) );
NAND2X1 NAND2X1_145 ( .A(cpuregs_5_[19]), .B(_5314__bF_buf1), .Y(_5334_) );
OAI21X1 OAI21X1_319 ( .A(_4793__bF_buf1), .B(_5314__bF_buf0), .C(_5334_), .Y(_205_) );
NAND2X1 NAND2X1_146 ( .A(cpuregs_5_[20]), .B(_5314__bF_buf7), .Y(_5335_) );
OAI21X1 OAI21X1_320 ( .A(_4806__bF_buf1), .B(_5314__bF_buf6), .C(_5335_), .Y(_206_) );
NAND2X1 NAND2X1_147 ( .A(cpuregs_5_[21]), .B(_5314__bF_buf5), .Y(_5336_) );
OAI21X1 OAI21X1_321 ( .A(_4816__bF_buf1), .B(_5314__bF_buf4), .C(_5336_), .Y(_207_) );
NAND2X1 NAND2X1_148 ( .A(cpuregs_5_[22]), .B(_5314__bF_buf3), .Y(_5337_) );
OAI21X1 OAI21X1_322 ( .A(_4824__bF_buf1), .B(_5314__bF_buf2), .C(_5337_), .Y(_208_) );
NAND2X1 NAND2X1_149 ( .A(cpuregs_5_[23]), .B(_5314__bF_buf1), .Y(_5338_) );
OAI21X1 OAI21X1_323 ( .A(_4833__bF_buf1), .B(_5314__bF_buf0), .C(_5338_), .Y(_209_) );
NAND2X1 NAND2X1_150 ( .A(cpuregs_5_[24]), .B(_5314__bF_buf7), .Y(_5339_) );
OAI21X1 OAI21X1_324 ( .A(_4845__bF_buf1), .B(_5314__bF_buf6), .C(_5339_), .Y(_210_) );
NAND2X1 NAND2X1_151 ( .A(cpuregs_5_[25]), .B(_5314__bF_buf5), .Y(_5340_) );
OAI21X1 OAI21X1_325 ( .A(_4854__bF_buf1), .B(_5314__bF_buf4), .C(_5340_), .Y(_211_) );
NAND2X1 NAND2X1_152 ( .A(cpuregs_5_[26]), .B(_5314__bF_buf3), .Y(_5341_) );
OAI21X1 OAI21X1_326 ( .A(_4863__bF_buf1), .B(_5314__bF_buf2), .C(_5341_), .Y(_212_) );
NAND2X1 NAND2X1_153 ( .A(cpuregs_5_[27]), .B(_5314__bF_buf1), .Y(_5342_) );
OAI21X1 OAI21X1_327 ( .A(_4871__bF_buf1), .B(_5314__bF_buf0), .C(_5342_), .Y(_213_) );
NAND2X1 NAND2X1_154 ( .A(cpuregs_5_[28]), .B(_5314__bF_buf7), .Y(_5343_) );
OAI21X1 OAI21X1_328 ( .A(_4884__bF_buf1), .B(_5314__bF_buf6), .C(_5343_), .Y(_214_) );
NAND2X1 NAND2X1_155 ( .A(cpuregs_5_[29]), .B(_5314__bF_buf5), .Y(_5344_) );
OAI21X1 OAI21X1_329 ( .A(_4893__bF_buf1), .B(_5314__bF_buf4), .C(_5344_), .Y(_215_) );
NAND2X1 NAND2X1_156 ( .A(cpuregs_5_[30]), .B(_5314__bF_buf3), .Y(_5345_) );
OAI21X1 OAI21X1_330 ( .A(_4901__bF_buf1), .B(_5314__bF_buf2), .C(_5345_), .Y(_216_) );
NAND2X1 NAND2X1_157 ( .A(cpuregs_5_[31]), .B(_5314__bF_buf1), .Y(_5346_) );
OAI21X1 OAI21X1_331 ( .A(_4910__bF_buf1), .B(_5314__bF_buf0), .C(_5346_), .Y(_217_) );
INVX1 INVX1_249 ( .A(decoded_rs2_4_bF_buf7_), .Y(_5347_) );
INVX1 INVX1_250 ( .A(decoded_rs2_3_bF_buf6_), .Y(_5348_) );
INVX1 INVX1_251 ( .A(decoded_rs2_1_bF_buf45_), .Y(_5349_) );
INVX1 INVX1_252 ( .A(cpuregs_12_[0]), .Y(_5350_) );
NAND2X1 NAND2X1_158 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_13_[0]), .Y(_5351_) );
OAI21X1 OAI21X1_332 ( .A(_5350_), .B(decoded_rs2_0_bF_buf77_), .C(_5351_), .Y(_5352_) );
INVX1 INVX1_253 ( .A(cpuregs_14_[0]), .Y(_5353_) );
NAND2X1 NAND2X1_159 ( .A(decoded_rs2_0_bF_buf76_), .B(cpuregs_15_[0]), .Y(_5354_) );
OAI21X1 OAI21X1_333 ( .A(_5353_), .B(decoded_rs2_0_bF_buf75_), .C(_5354_), .Y(_5355_) );
MUX2X1 MUX2X1_19 ( .A(_5352_), .B(_5355_), .S(_5349__bF_buf11), .Y(_5356_) );
NAND2X1 NAND2X1_160 ( .A(decoded_rs2_2_bF_buf8_), .B(_5356_), .Y(_5357_) );
INVX1 INVX1_254 ( .A(decoded_rs2_2_bF_buf7_), .Y(_5358_) );
INVX1 INVX1_255 ( .A(cpuregs_8_[0]), .Y(_5359_) );
NAND2X1 NAND2X1_161 ( .A(decoded_rs2_0_bF_buf74_), .B(cpuregs_9_[0]), .Y(_5360_) );
OAI21X1 OAI21X1_334 ( .A(_5359_), .B(decoded_rs2_0_bF_buf73_), .C(_5360_), .Y(_5361_) );
INVX1 INVX1_256 ( .A(decoded_rs2_0_bF_buf72_), .Y(_5362_) );
INVX1 INVX1_257 ( .A(cpuregs_11_[0]), .Y(_5363_) );
NAND2X1 NAND2X1_162 ( .A(cpuregs_10_[0]), .B(_5362__bF_buf14), .Y(_5364_) );
OAI21X1 OAI21X1_335 ( .A(_5362__bF_buf13), .B(_5363_), .C(_5364_), .Y(_5365_) );
MUX2X1 MUX2X1_20 ( .A(_5365_), .B(_5361_), .S(decoded_rs2_1_bF_buf44_), .Y(_5366_) );
AOI21X1 AOI21X1_28 ( .A(_5358__bF_buf12), .B(_5366_), .C(_5348__bF_buf5), .Y(_5367_) );
INVX1 INVX1_258 ( .A(cpuregs_4_[0]), .Y(_5368_) );
NAND2X1 NAND2X1_163 ( .A(cpuregs_5_[0]), .B(decoded_rs2_0_bF_buf71_), .Y(_5369_) );
OAI21X1 OAI21X1_336 ( .A(_5368_), .B(decoded_rs2_0_bF_buf70_), .C(_5369_), .Y(_5370_) );
NAND2X1 NAND2X1_164 ( .A(cpuregs_7_[0]), .B(decoded_rs2_0_bF_buf69_), .Y(_5371_) );
OAI21X1 OAI21X1_337 ( .A(_5269_), .B(decoded_rs2_0_bF_buf68_), .C(_5371_), .Y(_5372_) );
MUX2X1 MUX2X1_21 ( .A(_5372_), .B(_5370_), .S(decoded_rs2_1_bF_buf43_), .Y(_5373_) );
INVX1 INVX1_259 ( .A(cpuregs_0_[0]), .Y(_5374_) );
NAND2X1 NAND2X1_165 ( .A(cpuregs_1_[0]), .B(decoded_rs2_0_bF_buf67_), .Y(_5375_) );
OAI21X1 OAI21X1_338 ( .A(_5374_), .B(decoded_rs2_0_bF_buf66_), .C(_5375_), .Y(_5376_) );
INVX1 INVX1_260 ( .A(cpuregs_2_[0]), .Y(_5377_) );
NAND2X1 NAND2X1_166 ( .A(decoded_rs2_0_bF_buf65_), .B(cpuregs_3_[0]), .Y(_5378_) );
OAI21X1 OAI21X1_339 ( .A(_5377_), .B(decoded_rs2_0_bF_buf64_), .C(_5378_), .Y(_5379_) );
MUX2X1 MUX2X1_22 ( .A(_5376_), .B(_5379_), .S(_5349__bF_buf10), .Y(_5380_) );
MUX2X1 MUX2X1_23 ( .A(_5380_), .B(_5373_), .S(_5358__bF_buf11), .Y(_5381_) );
AOI22X1 AOI22X1_6 ( .A(_5348__bF_buf4), .B(_5381_), .C(_5367_), .D(_5357_), .Y(_5382_) );
NOR2X1 NOR2X1_236 ( .A(decoded_rs2_0_bF_buf63_), .B(decoded_rs2_1_bF_buf42_), .Y(_5383_) );
INVX1 INVX1_261 ( .A(_5383_), .Y(_5384_) );
NAND3X1 NAND3X1_21 ( .A(_5358__bF_buf10), .B(_5348__bF_buf3), .C(_5347_), .Y(_5385_) );
INVX1 INVX1_262 ( .A(cpuregs_26_[0]), .Y(_5386_) );
OAI21X1 OAI21X1_340 ( .A(_5386_), .B(decoded_rs2_0_bF_buf62_), .C(decoded_rs2_1_bF_buf41_), .Y(_5387_) );
AOI21X1 AOI21X1_29 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_27_[0]), .C(_5387_), .Y(_5388_) );
AND2X2 AND2X2_18 ( .A(decoded_rs2_0_bF_buf60_), .B(cpuregs_25_[0]), .Y(_5389_) );
INVX1 INVX1_263 ( .A(cpuregs_24_[0]), .Y(_5390_) );
OAI21X1 OAI21X1_341 ( .A(_5390_), .B(decoded_rs2_0_bF_buf59_), .C(_5349__bF_buf9), .Y(_5391_) );
OAI21X1 OAI21X1_342 ( .A(_5391_), .B(_5389_), .C(_5358__bF_buf9), .Y(_5392_) );
INVX1 INVX1_264 ( .A(cpuregs_30_[0]), .Y(_5393_) );
OAI21X1 OAI21X1_343 ( .A(_5393_), .B(decoded_rs2_0_bF_buf58_), .C(decoded_rs2_1_bF_buf40_), .Y(_5394_) );
AOI21X1 AOI21X1_30 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_31_[0]), .C(_5394_), .Y(_5395_) );
AND2X2 AND2X2_19 ( .A(_5362__bF_buf12), .B(cpuregs_28_[0]), .Y(_5396_) );
INVX1 INVX1_265 ( .A(cpuregs_29_[0]), .Y(_5397_) );
OAI21X1 OAI21X1_344 ( .A(_5362__bF_buf11), .B(_5397_), .C(_5349__bF_buf8), .Y(_5398_) );
OAI21X1 OAI21X1_345 ( .A(_5398_), .B(_5396_), .C(decoded_rs2_2_bF_buf6_), .Y(_5399_) );
OAI22X1 OAI22X1_4 ( .A(_5392_), .B(_5388_), .C(_5399_), .D(_5395_), .Y(_5400_) );
INVX1 INVX1_266 ( .A(cpuregs_16_[0]), .Y(_5401_) );
NAND2X1 NAND2X1_167 ( .A(decoded_rs2_0_bF_buf56_), .B(cpuregs_17_[0]), .Y(_5402_) );
OAI21X1 OAI21X1_346 ( .A(_5401_), .B(decoded_rs2_0_bF_buf55_), .C(_5402_), .Y(_5403_) );
INVX1 INVX1_267 ( .A(cpuregs_18_[0]), .Y(_5404_) );
NAND2X1 NAND2X1_168 ( .A(decoded_rs2_0_bF_buf54_), .B(cpuregs_19_[0]), .Y(_5405_) );
OAI21X1 OAI21X1_347 ( .A(_5404_), .B(decoded_rs2_0_bF_buf53_), .C(_5405_), .Y(_5406_) );
MUX2X1 MUX2X1_24 ( .A(_5403_), .B(_5406_), .S(_5349__bF_buf7), .Y(_5407_) );
INVX1 INVX1_268 ( .A(cpuregs_20_[0]), .Y(_5408_) );
NAND2X1 NAND2X1_169 ( .A(decoded_rs2_0_bF_buf52_), .B(cpuregs_21_[0]), .Y(_5409_) );
OAI21X1 OAI21X1_348 ( .A(_5408_), .B(decoded_rs2_0_bF_buf51_), .C(_5409_), .Y(_5410_) );
INVX1 INVX1_269 ( .A(cpuregs_22_[0]), .Y(_5411_) );
NAND2X1 NAND2X1_170 ( .A(decoded_rs2_0_bF_buf50_), .B(cpuregs_23_[0]), .Y(_5412_) );
OAI21X1 OAI21X1_349 ( .A(_5411_), .B(decoded_rs2_0_bF_buf49_), .C(_5412_), .Y(_5413_) );
MUX2X1 MUX2X1_25 ( .A(_5410_), .B(_5413_), .S(_5349__bF_buf6), .Y(_5414_) );
MUX2X1 MUX2X1_26 ( .A(_5414_), .B(_5407_), .S(decoded_rs2_2_bF_buf5_), .Y(_5415_) );
MUX2X1 MUX2X1_27 ( .A(_5400_), .B(_5415_), .S(decoded_rs2_3_bF_buf5_), .Y(_5416_) );
NAND2X1 NAND2X1_171 ( .A(decoded_rs2_4_bF_buf6_), .B(_5416_), .Y(_5417_) );
OAI21X1 OAI21X1_350 ( .A(_5384_), .B(_5385_), .C(_5417_), .Y(_5418_) );
AOI21X1 AOI21X1_31 ( .A(_5347_), .B(_5382_), .C(_5418_), .Y(_5419_) );
NAND2X1 NAND2X1_172 ( .A(is_slli_srli_srai), .B(_5362__bF_buf10), .Y(_5420_) );
OAI21X1 OAI21X1_351 ( .A(_5419_), .B(is_slli_srli_srai), .C(_5420_), .Y(_5421_) );
AND2X2 AND2X2_20 ( .A(_4580__bF_buf3), .B(reg_sh_0_), .Y(_5422_) );
OAI21X1 OAI21X1_352 ( .A(_5422_), .B(_4581_), .C(cpu_state_4_), .Y(_5423_) );
OAI21X1 OAI21X1_353 ( .A(_5421_), .B(cpu_state_4_), .C(_5423_), .Y(_85__0_) );
INVX1 INVX1_270 ( .A(cpuregs_12_[1]), .Y(_5424_) );
NAND2X1 NAND2X1_173 ( .A(decoded_rs2_0_bF_buf48_), .B(cpuregs_13_[1]), .Y(_5425_) );
OAI21X1 OAI21X1_354 ( .A(_5424_), .B(decoded_rs2_0_bF_buf47_), .C(_5425_), .Y(_5426_) );
INVX1 INVX1_271 ( .A(cpuregs_14_[1]), .Y(_5427_) );
NAND2X1 NAND2X1_174 ( .A(decoded_rs2_0_bF_buf46_), .B(cpuregs_15_[1]), .Y(_5428_) );
OAI21X1 OAI21X1_355 ( .A(_5427_), .B(decoded_rs2_0_bF_buf45_), .C(_5428_), .Y(_5429_) );
MUX2X1 MUX2X1_28 ( .A(_5429_), .B(_5426_), .S(decoded_rs2_1_bF_buf39_), .Y(_5430_) );
NAND2X1 NAND2X1_175 ( .A(decoded_rs2_2_bF_buf4_), .B(_5430_), .Y(_5431_) );
INVX1 INVX1_272 ( .A(cpuregs_8_[1]), .Y(_5432_) );
NAND2X1 NAND2X1_176 ( .A(decoded_rs2_0_bF_buf44_), .B(cpuregs_9_[1]), .Y(_5433_) );
OAI21X1 OAI21X1_356 ( .A(_5432_), .B(decoded_rs2_0_bF_buf43_), .C(_5433_), .Y(_5434_) );
INVX1 INVX1_273 ( .A(cpuregs_10_[1]), .Y(_5435_) );
NAND2X1 NAND2X1_177 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_11_[1]), .Y(_5436_) );
OAI21X1 OAI21X1_357 ( .A(_5435_), .B(decoded_rs2_0_bF_buf41_), .C(_5436_), .Y(_5437_) );
MUX2X1 MUX2X1_29 ( .A(_5437_), .B(_5434_), .S(decoded_rs2_1_bF_buf38_), .Y(_5438_) );
AOI21X1 AOI21X1_32 ( .A(_5358__bF_buf8), .B(_5438_), .C(_5348__bF_buf2), .Y(_5439_) );
INVX1 INVX1_274 ( .A(cpuregs_4_[1]), .Y(_5440_) );
NAND2X1 NAND2X1_178 ( .A(cpuregs_5_[1]), .B(decoded_rs2_0_bF_buf40_), .Y(_5441_) );
OAI21X1 OAI21X1_358 ( .A(_5440_), .B(decoded_rs2_0_bF_buf39_), .C(_5441_), .Y(_5442_) );
NAND2X1 NAND2X1_179 ( .A(cpuregs_7_[1]), .B(decoded_rs2_0_bF_buf38_), .Y(_5443_) );
OAI21X1 OAI21X1_359 ( .A(_5275_), .B(decoded_rs2_0_bF_buf37_), .C(_5443_), .Y(_5444_) );
MUX2X1 MUX2X1_30 ( .A(_5444_), .B(_5442_), .S(decoded_rs2_1_bF_buf37_), .Y(_5445_) );
NOR2X1 NOR2X1_237 ( .A(decoded_rs2_0_bF_buf36_), .B(cpuregs_0_[1]), .Y(_5446_) );
OAI21X1 OAI21X1_360 ( .A(_5362__bF_buf9), .B(cpuregs_1_[1]), .C(_5349__bF_buf5), .Y(_5447_) );
NOR2X1 NOR2X1_238 ( .A(_5446_), .B(_5447_), .Y(_5448_) );
INVX1 INVX1_275 ( .A(cpuregs_3_[1]), .Y(_5449_) );
OAI21X1 OAI21X1_361 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_2_[1]), .C(decoded_rs2_1_bF_buf36_), .Y(_5450_) );
AOI21X1 AOI21X1_33 ( .A(decoded_rs2_0_bF_buf34_), .B(_5449_), .C(_5450_), .Y(_5451_) );
OAI21X1 OAI21X1_362 ( .A(_5448_), .B(_5451_), .C(_5358__bF_buf7), .Y(_5452_) );
OAI21X1 OAI21X1_363 ( .A(_5358__bF_buf6), .B(_5445_), .C(_5452_), .Y(_5453_) );
AOI22X1 AOI22X1_7 ( .A(_5431_), .B(_5439_), .C(_5453_), .D(_5348__bF_buf1), .Y(_5454_) );
INVX1 INVX1_276 ( .A(cpuregs_26_[1]), .Y(_5455_) );
OAI21X1 OAI21X1_364 ( .A(_5455_), .B(decoded_rs2_0_bF_buf33_), .C(decoded_rs2_1_bF_buf35_), .Y(_5456_) );
AOI21X1 AOI21X1_34 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_27_[1]), .C(_5456_), .Y(_5457_) );
AND2X2 AND2X2_21 ( .A(decoded_rs2_0_bF_buf31_), .B(cpuregs_25_[1]), .Y(_5458_) );
INVX1 INVX1_277 ( .A(cpuregs_24_[1]), .Y(_5459_) );
OAI21X1 OAI21X1_365 ( .A(_5459_), .B(decoded_rs2_0_bF_buf30_), .C(_5349__bF_buf4), .Y(_5460_) );
OAI21X1 OAI21X1_366 ( .A(_5460_), .B(_5458_), .C(_5358__bF_buf5), .Y(_5461_) );
INVX1 INVX1_278 ( .A(cpuregs_28_[1]), .Y(_5462_) );
NAND2X1 NAND2X1_180 ( .A(decoded_rs2_0_bF_buf29_), .B(cpuregs_29_[1]), .Y(_5463_) );
OAI21X1 OAI21X1_367 ( .A(_5462_), .B(decoded_rs2_0_bF_buf28_), .C(_5463_), .Y(_5464_) );
INVX1 INVX1_279 ( .A(cpuregs_30_[1]), .Y(_5465_) );
NAND2X1 NAND2X1_181 ( .A(decoded_rs2_0_bF_buf27_), .B(cpuregs_31_[1]), .Y(_5466_) );
OAI21X1 OAI21X1_368 ( .A(_5465_), .B(decoded_rs2_0_bF_buf26_), .C(_5466_), .Y(_5467_) );
MUX2X1 MUX2X1_31 ( .A(_5467_), .B(_5464_), .S(decoded_rs2_1_bF_buf34_), .Y(_5468_) );
OAI22X1 OAI22X1_5 ( .A(_5461_), .B(_5457_), .C(_5468_), .D(_5358__bF_buf4), .Y(_5469_) );
INVX1 INVX1_280 ( .A(cpuregs_16_[1]), .Y(_5470_) );
NAND2X1 NAND2X1_182 ( .A(decoded_rs2_0_bF_buf25_), .B(cpuregs_17_[1]), .Y(_5471_) );
OAI21X1 OAI21X1_369 ( .A(_5470_), .B(decoded_rs2_0_bF_buf24_), .C(_5471_), .Y(_5472_) );
INVX1 INVX1_281 ( .A(cpuregs_18_[1]), .Y(_5473_) );
NAND2X1 NAND2X1_183 ( .A(decoded_rs2_0_bF_buf23_), .B(cpuregs_19_[1]), .Y(_5474_) );
OAI21X1 OAI21X1_370 ( .A(_5473_), .B(decoded_rs2_0_bF_buf22_), .C(_5474_), .Y(_5475_) );
MUX2X1 MUX2X1_32 ( .A(_5475_), .B(_5472_), .S(decoded_rs2_1_bF_buf33_), .Y(_5476_) );
INVX1 INVX1_282 ( .A(cpuregs_20_[1]), .Y(_5477_) );
NAND2X1 NAND2X1_184 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_21_[1]), .Y(_5478_) );
OAI21X1 OAI21X1_371 ( .A(_5477_), .B(decoded_rs2_0_bF_buf20_), .C(_5478_), .Y(_5479_) );
INVX1 INVX1_283 ( .A(cpuregs_23_[1]), .Y(_5480_) );
NAND2X1 NAND2X1_185 ( .A(cpuregs_22_[1]), .B(_5362__bF_buf8), .Y(_5481_) );
OAI21X1 OAI21X1_372 ( .A(_5362__bF_buf7), .B(_5480_), .C(_5481_), .Y(_5482_) );
MUX2X1 MUX2X1_33 ( .A(_5482_), .B(_5479_), .S(decoded_rs2_1_bF_buf32_), .Y(_5483_) );
MUX2X1 MUX2X1_34 ( .A(_5483_), .B(_5476_), .S(decoded_rs2_2_bF_buf3_), .Y(_5484_) );
MUX2X1 MUX2X1_35 ( .A(_5484_), .B(_5469_), .S(_5348__bF_buf0), .Y(_5485_) );
NAND2X1 NAND2X1_186 ( .A(decoded_rs2_4_bF_buf5_), .B(_5485_), .Y(_5486_) );
OAI21X1 OAI21X1_373 ( .A(_5384_), .B(_5385_), .C(_5486_), .Y(_5487_) );
AOI21X1 AOI21X1_35 ( .A(_5347_), .B(_5454_), .C(_5487_), .Y(_5488_) );
NOR2X1 NOR2X1_239 ( .A(is_slli_srli_srai), .B(_5488_), .Y(_5489_) );
OAI21X1 OAI21X1_374 ( .A(_4564_), .B(decoded_rs2_1_bF_buf31_), .C(_4575__bF_buf2), .Y(_5490_) );
NOR2X1 NOR2X1_240 ( .A(_4576_), .B(_4581_), .Y(_5491_) );
OAI21X1 OAI21X1_375 ( .A(_4583_), .B(_5491_), .C(cpu_state_4_), .Y(_5492_) );
OAI21X1 OAI21X1_376 ( .A(_5489_), .B(_5490_), .C(_5492_), .Y(_85__1_) );
INVX1 INVX1_284 ( .A(cpuregs_12_[2]), .Y(_5493_) );
NAND2X1 NAND2X1_187 ( .A(decoded_rs2_0_bF_buf19_), .B(cpuregs_13_[2]), .Y(_5494_) );
OAI21X1 OAI21X1_377 ( .A(_5493_), .B(decoded_rs2_0_bF_buf18_), .C(_5494_), .Y(_5495_) );
INVX1 INVX1_285 ( .A(cpuregs_14_[2]), .Y(_5496_) );
NAND2X1 NAND2X1_188 ( .A(decoded_rs2_0_bF_buf17_), .B(cpuregs_15_[2]), .Y(_5497_) );
OAI21X1 OAI21X1_378 ( .A(_5496_), .B(decoded_rs2_0_bF_buf16_), .C(_5497_), .Y(_5498_) );
MUX2X1 MUX2X1_36 ( .A(_5498_), .B(_5495_), .S(decoded_rs2_1_bF_buf30_), .Y(_5499_) );
NAND2X1 NAND2X1_189 ( .A(decoded_rs2_2_bF_buf2_), .B(_5499_), .Y(_5500_) );
INVX1 INVX1_286 ( .A(cpuregs_8_[2]), .Y(_5501_) );
NAND2X1 NAND2X1_190 ( .A(decoded_rs2_0_bF_buf15_), .B(cpuregs_9_[2]), .Y(_5502_) );
OAI21X1 OAI21X1_379 ( .A(_5501_), .B(decoded_rs2_0_bF_buf14_), .C(_5502_), .Y(_5503_) );
INVX1 INVX1_287 ( .A(cpuregs_10_[2]), .Y(_5504_) );
NAND2X1 NAND2X1_191 ( .A(decoded_rs2_0_bF_buf13_), .B(cpuregs_11_[2]), .Y(_5505_) );
OAI21X1 OAI21X1_380 ( .A(_5504_), .B(decoded_rs2_0_bF_buf12_), .C(_5505_), .Y(_5506_) );
MUX2X1 MUX2X1_37 ( .A(_5506_), .B(_5503_), .S(decoded_rs2_1_bF_buf29_), .Y(_5507_) );
AOI21X1 AOI21X1_36 ( .A(_5358__bF_buf3), .B(_5507_), .C(_5348__bF_buf5), .Y(_5508_) );
INVX1 INVX1_288 ( .A(cpuregs_4_[2]), .Y(_5509_) );
NAND2X1 NAND2X1_192 ( .A(cpuregs_5_[2]), .B(decoded_rs2_0_bF_buf11_), .Y(_5510_) );
OAI21X1 OAI21X1_381 ( .A(_5509_), .B(decoded_rs2_0_bF_buf10_), .C(_5510_), .Y(_5511_) );
NAND2X1 NAND2X1_193 ( .A(cpuregs_7_[2]), .B(decoded_rs2_0_bF_buf9_), .Y(_5512_) );
OAI21X1 OAI21X1_382 ( .A(_5276_), .B(decoded_rs2_0_bF_buf8_), .C(_5512_), .Y(_5513_) );
MUX2X1 MUX2X1_38 ( .A(_5513_), .B(_5511_), .S(decoded_rs2_1_bF_buf28_), .Y(_5514_) );
NOR2X1 NOR2X1_241 ( .A(decoded_rs2_0_bF_buf7_), .B(cpuregs_0_[2]), .Y(_5515_) );
OAI21X1 OAI21X1_383 ( .A(_5362__bF_buf6), .B(cpuregs_1_[2]), .C(_5349__bF_buf3), .Y(_5516_) );
NOR2X1 NOR2X1_242 ( .A(_5515_), .B(_5516_), .Y(_5517_) );
INVX1 INVX1_289 ( .A(cpuregs_3_[2]), .Y(_5518_) );
OAI21X1 OAI21X1_384 ( .A(decoded_rs2_0_bF_buf6_), .B(cpuregs_2_[2]), .C(decoded_rs2_1_bF_buf27_), .Y(_5519_) );
AOI21X1 AOI21X1_37 ( .A(decoded_rs2_0_bF_buf5_), .B(_5518_), .C(_5519_), .Y(_5520_) );
OAI21X1 OAI21X1_385 ( .A(_5517_), .B(_5520_), .C(_5358__bF_buf2), .Y(_5521_) );
OAI21X1 OAI21X1_386 ( .A(_5358__bF_buf1), .B(_5514_), .C(_5521_), .Y(_5522_) );
AOI22X1 AOI22X1_8 ( .A(_5500_), .B(_5508_), .C(_5522_), .D(_5348__bF_buf4), .Y(_5523_) );
INVX1 INVX1_290 ( .A(cpuregs_31_[2]), .Y(_5524_) );
OAI21X1 OAI21X1_387 ( .A(_5358__bF_buf0), .B(_5524_), .C(decoded_rs2_0_bF_buf4_), .Y(_5525_) );
AOI21X1 AOI21X1_38 ( .A(_5358__bF_buf12), .B(cpuregs_27_[2]), .C(_5525_), .Y(_5526_) );
INVX1 INVX1_291 ( .A(cpuregs_26_[2]), .Y(_5527_) );
NOR2X1 NOR2X1_243 ( .A(decoded_rs2_2_bF_buf1_), .B(_5527_), .Y(_5528_) );
INVX1 INVX1_292 ( .A(cpuregs_30_[2]), .Y(_5529_) );
OAI21X1 OAI21X1_388 ( .A(_5358__bF_buf11), .B(_5529_), .C(_5362__bF_buf5), .Y(_5530_) );
OAI21X1 OAI21X1_389 ( .A(_5530_), .B(_5528_), .C(decoded_rs2_1_bF_buf26_), .Y(_5531_) );
INVX1 INVX1_293 ( .A(cpuregs_29_[2]), .Y(_5532_) );
OAI21X1 OAI21X1_390 ( .A(_5358__bF_buf10), .B(_5532_), .C(decoded_rs2_0_bF_buf3_), .Y(_5533_) );
AOI21X1 AOI21X1_39 ( .A(_5358__bF_buf9), .B(cpuregs_25_[2]), .C(_5533_), .Y(_5534_) );
INVX1 INVX1_294 ( .A(cpuregs_24_[2]), .Y(_5535_) );
NOR2X1 NOR2X1_244 ( .A(decoded_rs2_2_bF_buf0_), .B(_5535_), .Y(_5536_) );
INVX1 INVX1_295 ( .A(cpuregs_28_[2]), .Y(_5537_) );
OAI21X1 OAI21X1_391 ( .A(_5358__bF_buf8), .B(_5537_), .C(_5362__bF_buf4), .Y(_5538_) );
OAI21X1 OAI21X1_392 ( .A(_5538_), .B(_5536_), .C(_5349__bF_buf2), .Y(_5539_) );
OAI22X1 OAI22X1_6 ( .A(_5531_), .B(_5526_), .C(_5534_), .D(_5539_), .Y(_5540_) );
INVX1 INVX1_296 ( .A(cpuregs_16_[2]), .Y(_5541_) );
NAND2X1 NAND2X1_194 ( .A(decoded_rs2_0_bF_buf2_), .B(cpuregs_17_[2]), .Y(_5542_) );
OAI21X1 OAI21X1_393 ( .A(_5541_), .B(decoded_rs2_0_bF_buf1_), .C(_5542_), .Y(_5543_) );
INVX1 INVX1_297 ( .A(cpuregs_18_[2]), .Y(_5544_) );
NAND2X1 NAND2X1_195 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_19_[2]), .Y(_5545_) );
OAI21X1 OAI21X1_394 ( .A(_5544_), .B(decoded_rs2_0_bF_buf78_), .C(_5545_), .Y(_5546_) );
MUX2X1 MUX2X1_39 ( .A(_5546_), .B(_5543_), .S(decoded_rs2_1_bF_buf25_), .Y(_5547_) );
NAND2X1 NAND2X1_196 ( .A(_5358__bF_buf7), .B(_5547_), .Y(_5548_) );
INVX1 INVX1_298 ( .A(cpuregs_20_[2]), .Y(_5549_) );
NAND2X1 NAND2X1_197 ( .A(decoded_rs2_0_bF_buf77_), .B(cpuregs_21_[2]), .Y(_5550_) );
OAI21X1 OAI21X1_395 ( .A(_5549_), .B(decoded_rs2_0_bF_buf76_), .C(_5550_), .Y(_5551_) );
INVX1 INVX1_299 ( .A(cpuregs_22_[2]), .Y(_5552_) );
NAND2X1 NAND2X1_198 ( .A(decoded_rs2_0_bF_buf75_), .B(cpuregs_23_[2]), .Y(_5553_) );
OAI21X1 OAI21X1_396 ( .A(_5552_), .B(decoded_rs2_0_bF_buf74_), .C(_5553_), .Y(_5554_) );
MUX2X1 MUX2X1_40 ( .A(_5554_), .B(_5551_), .S(decoded_rs2_1_bF_buf24_), .Y(_5555_) );
AOI21X1 AOI21X1_40 ( .A(decoded_rs2_2_bF_buf8_), .B(_5555_), .C(decoded_rs2_3_bF_buf4_), .Y(_5556_) );
AOI22X1 AOI22X1_9 ( .A(_5548_), .B(_5556_), .C(_5540_), .D(decoded_rs2_3_bF_buf3_), .Y(_5557_) );
NAND2X1 NAND2X1_199 ( .A(decoded_rs2_4_bF_buf4_), .B(_5557_), .Y(_5558_) );
OAI21X1 OAI21X1_397 ( .A(_5384_), .B(_5385_), .C(_5558_), .Y(_5559_) );
AOI21X1 AOI21X1_41 ( .A(_5347_), .B(_5523_), .C(_5559_), .Y(_5560_) );
NOR2X1 NOR2X1_245 ( .A(is_slli_srli_srai), .B(_5560_), .Y(_5561_) );
OAI21X1 OAI21X1_398 ( .A(_4564_), .B(decoded_rs2_2_bF_buf7_), .C(_4575__bF_buf1), .Y(_5562_) );
OAI21X1 OAI21X1_399 ( .A(reg_sh_2_), .B(_4579__bF_buf3), .C(_4582_), .Y(_5563_) );
NAND2X1 NAND2X1_200 ( .A(cpu_state_4_), .B(_5563_), .Y(_5564_) );
OAI21X1 OAI21X1_400 ( .A(_5561_), .B(_5562_), .C(_5564_), .Y(_85__2_) );
INVX1 INVX1_300 ( .A(cpuregs_12_[3]), .Y(_5565_) );
NAND2X1 NAND2X1_201 ( .A(decoded_rs2_0_bF_buf73_), .B(cpuregs_13_[3]), .Y(_5566_) );
OAI21X1 OAI21X1_401 ( .A(_5565_), .B(decoded_rs2_0_bF_buf72_), .C(_5566_), .Y(_5567_) );
INVX1 INVX1_301 ( .A(cpuregs_14_[3]), .Y(_5568_) );
NAND2X1 NAND2X1_202 ( .A(decoded_rs2_0_bF_buf71_), .B(cpuregs_15_[3]), .Y(_5569_) );
OAI21X1 OAI21X1_402 ( .A(_5568_), .B(decoded_rs2_0_bF_buf70_), .C(_5569_), .Y(_5570_) );
MUX2X1 MUX2X1_41 ( .A(_5570_), .B(_5567_), .S(decoded_rs2_1_bF_buf23_), .Y(_5571_) );
NAND2X1 NAND2X1_203 ( .A(decoded_rs2_2_bF_buf6_), .B(_5571_), .Y(_5572_) );
INVX1 INVX1_302 ( .A(cpuregs_8_[3]), .Y(_5573_) );
NAND2X1 NAND2X1_204 ( .A(decoded_rs2_0_bF_buf69_), .B(cpuregs_9_[3]), .Y(_5574_) );
OAI21X1 OAI21X1_403 ( .A(_5573_), .B(decoded_rs2_0_bF_buf68_), .C(_5574_), .Y(_5575_) );
INVX1 INVX1_303 ( .A(cpuregs_10_[3]), .Y(_5576_) );
NAND2X1 NAND2X1_205 ( .A(decoded_rs2_0_bF_buf67_), .B(cpuregs_11_[3]), .Y(_5577_) );
OAI21X1 OAI21X1_404 ( .A(_5576_), .B(decoded_rs2_0_bF_buf66_), .C(_5577_), .Y(_5578_) );
MUX2X1 MUX2X1_42 ( .A(_5578_), .B(_5575_), .S(decoded_rs2_1_bF_buf22_), .Y(_5579_) );
AOI21X1 AOI21X1_42 ( .A(_5358__bF_buf6), .B(_5579_), .C(_5348__bF_buf3), .Y(_5580_) );
INVX1 INVX1_304 ( .A(cpuregs_4_[3]), .Y(_5581_) );
NAND2X1 NAND2X1_206 ( .A(cpuregs_5_[3]), .B(decoded_rs2_0_bF_buf65_), .Y(_5582_) );
OAI21X1 OAI21X1_405 ( .A(_5581_), .B(decoded_rs2_0_bF_buf64_), .C(_5582_), .Y(_5583_) );
NAND2X1 NAND2X1_207 ( .A(cpuregs_7_[3]), .B(decoded_rs2_0_bF_buf63_), .Y(_5584_) );
OAI21X1 OAI21X1_406 ( .A(_5277_), .B(decoded_rs2_0_bF_buf62_), .C(_5584_), .Y(_5585_) );
MUX2X1 MUX2X1_43 ( .A(_5585_), .B(_5583_), .S(decoded_rs2_1_bF_buf21_), .Y(_5586_) );
NOR2X1 NOR2X1_246 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_0_[3]), .Y(_5587_) );
OAI21X1 OAI21X1_407 ( .A(_5362__bF_buf3), .B(cpuregs_1_[3]), .C(_5349__bF_buf1), .Y(_5588_) );
NOR2X1 NOR2X1_247 ( .A(_5587_), .B(_5588_), .Y(_5589_) );
INVX1 INVX1_305 ( .A(cpuregs_3_[3]), .Y(_5590_) );
OAI21X1 OAI21X1_408 ( .A(decoded_rs2_0_bF_buf60_), .B(cpuregs_2_[3]), .C(decoded_rs2_1_bF_buf20_), .Y(_5591_) );
AOI21X1 AOI21X1_43 ( .A(decoded_rs2_0_bF_buf59_), .B(_5590_), .C(_5591_), .Y(_5592_) );
OAI21X1 OAI21X1_409 ( .A(_5589_), .B(_5592_), .C(_5358__bF_buf5), .Y(_5593_) );
OAI21X1 OAI21X1_410 ( .A(_5358__bF_buf4), .B(_5586_), .C(_5593_), .Y(_5594_) );
AOI22X1 AOI22X1_10 ( .A(_5572_), .B(_5580_), .C(_5594_), .D(_5348__bF_buf2), .Y(_5595_) );
NOR2X1 NOR2X1_248 ( .A(decoded_rs2_0_bF_buf58_), .B(cpuregs_24_[3]), .Y(_5596_) );
OAI21X1 OAI21X1_411 ( .A(_5362__bF_buf2), .B(cpuregs_25_[3]), .C(_5349__bF_buf0), .Y(_5597_) );
NOR2X1 NOR2X1_249 ( .A(_5596_), .B(_5597_), .Y(_5598_) );
INVX1 INVX1_306 ( .A(cpuregs_27_[3]), .Y(_5599_) );
OAI21X1 OAI21X1_412 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_26_[3]), .C(decoded_rs2_1_bF_buf19_), .Y(_5600_) );
AOI21X1 AOI21X1_44 ( .A(decoded_rs2_0_bF_buf56_), .B(_5599_), .C(_5600_), .Y(_5601_) );
OAI21X1 OAI21X1_413 ( .A(_5598_), .B(_5601_), .C(_5358__bF_buf3), .Y(_5602_) );
INVX1 INVX1_307 ( .A(cpuregs_28_[3]), .Y(_5603_) );
OAI21X1 OAI21X1_414 ( .A(_5362__bF_buf1), .B(cpuregs_29_[3]), .C(_5349__bF_buf11), .Y(_5604_) );
AOI21X1 AOI21X1_45 ( .A(_5362__bF_buf0), .B(_5603_), .C(_5604_), .Y(_5605_) );
INVX1 INVX1_308 ( .A(cpuregs_31_[3]), .Y(_5606_) );
OAI21X1 OAI21X1_415 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_30_[3]), .C(decoded_rs2_1_bF_buf18_), .Y(_5607_) );
AOI21X1 AOI21X1_46 ( .A(decoded_rs2_0_bF_buf54_), .B(_5606_), .C(_5607_), .Y(_5608_) );
OAI21X1 OAI21X1_416 ( .A(_5605_), .B(_5608_), .C(decoded_rs2_2_bF_buf5_), .Y(_5609_) );
AOI21X1 AOI21X1_47 ( .A(_5602_), .B(_5609_), .C(_5348__bF_buf1), .Y(_5610_) );
INVX1 INVX1_309 ( .A(cpuregs_16_[3]), .Y(_5611_) );
NAND2X1 NAND2X1_208 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_17_[3]), .Y(_5612_) );
OAI21X1 OAI21X1_417 ( .A(_5611_), .B(decoded_rs2_0_bF_buf52_), .C(_5612_), .Y(_5613_) );
INVX1 INVX1_310 ( .A(cpuregs_18_[3]), .Y(_5614_) );
NAND2X1 NAND2X1_209 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_19_[3]), .Y(_5615_) );
OAI21X1 OAI21X1_418 ( .A(_5614_), .B(decoded_rs2_0_bF_buf50_), .C(_5615_), .Y(_5616_) );
MUX2X1 MUX2X1_44 ( .A(_5616_), .B(_5613_), .S(decoded_rs2_1_bF_buf17_), .Y(_5617_) );
INVX1 INVX1_311 ( .A(cpuregs_20_[3]), .Y(_5618_) );
NAND2X1 NAND2X1_210 ( .A(decoded_rs2_0_bF_buf49_), .B(cpuregs_21_[3]), .Y(_5619_) );
OAI21X1 OAI21X1_419 ( .A(_5618_), .B(decoded_rs2_0_bF_buf48_), .C(_5619_), .Y(_5620_) );
INVX1 INVX1_312 ( .A(cpuregs_23_[3]), .Y(_5621_) );
NAND2X1 NAND2X1_211 ( .A(cpuregs_22_[3]), .B(_5362__bF_buf14), .Y(_5622_) );
OAI21X1 OAI21X1_420 ( .A(_5362__bF_buf13), .B(_5621_), .C(_5622_), .Y(_5623_) );
MUX2X1 MUX2X1_45 ( .A(_5623_), .B(_5620_), .S(decoded_rs2_1_bF_buf16_), .Y(_5624_) );
MUX2X1 MUX2X1_46 ( .A(_5624_), .B(_5617_), .S(decoded_rs2_2_bF_buf4_), .Y(_5625_) );
AOI21X1 AOI21X1_48 ( .A(_5348__bF_buf0), .B(_5625_), .C(_5610_), .Y(_5626_) );
NAND2X1 NAND2X1_212 ( .A(decoded_rs2_4_bF_buf3_), .B(_5626_), .Y(_5627_) );
OAI21X1 OAI21X1_421 ( .A(_5384_), .B(_5385_), .C(_5627_), .Y(_5628_) );
AOI21X1 AOI21X1_49 ( .A(_5347_), .B(_5595_), .C(_5628_), .Y(_5629_) );
NOR2X1 NOR2X1_250 ( .A(is_slli_srli_srai), .B(_5629_), .Y(_5630_) );
OAI21X1 OAI21X1_422 ( .A(_4564_), .B(decoded_rs2_3_bF_buf2_), .C(_4575__bF_buf0), .Y(_5631_) );
INVX1 INVX1_313 ( .A(reg_sh_4_), .Y(_5632_) );
NAND2X1 NAND2X1_213 ( .A(reg_sh_3_), .B(reg_sh_2_), .Y(_5633_) );
OAI21X1 OAI21X1_423 ( .A(_4578_), .B(_5632_), .C(_5633_), .Y(_5634_) );
OAI21X1 OAI21X1_424 ( .A(_4583_), .B(_5634_), .C(cpu_state_4_), .Y(_5635_) );
OAI21X1 OAI21X1_425 ( .A(_5630_), .B(_5631_), .C(_5635_), .Y(_85__3_) );
INVX1 INVX1_314 ( .A(cpuregs_12_[4]), .Y(_5636_) );
NAND2X1 NAND2X1_214 ( .A(decoded_rs2_0_bF_buf47_), .B(cpuregs_13_[4]), .Y(_5637_) );
OAI21X1 OAI21X1_426 ( .A(_5636_), .B(decoded_rs2_0_bF_buf46_), .C(_5637_), .Y(_5638_) );
INVX1 INVX1_315 ( .A(cpuregs_14_[4]), .Y(_5639_) );
NAND2X1 NAND2X1_215 ( .A(decoded_rs2_0_bF_buf45_), .B(cpuregs_15_[4]), .Y(_5640_) );
OAI21X1 OAI21X1_427 ( .A(_5639_), .B(decoded_rs2_0_bF_buf44_), .C(_5640_), .Y(_5641_) );
MUX2X1 MUX2X1_47 ( .A(_5641_), .B(_5638_), .S(decoded_rs2_1_bF_buf15_), .Y(_5642_) );
NAND2X1 NAND2X1_216 ( .A(decoded_rs2_2_bF_buf3_), .B(_5642_), .Y(_5643_) );
INVX1 INVX1_316 ( .A(cpuregs_8_[4]), .Y(_5644_) );
NAND2X1 NAND2X1_217 ( .A(decoded_rs2_0_bF_buf43_), .B(cpuregs_9_[4]), .Y(_5645_) );
OAI21X1 OAI21X1_428 ( .A(_5644_), .B(decoded_rs2_0_bF_buf42_), .C(_5645_), .Y(_5646_) );
INVX1 INVX1_317 ( .A(cpuregs_10_[4]), .Y(_5647_) );
NAND2X1 NAND2X1_218 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_11_[4]), .Y(_5648_) );
OAI21X1 OAI21X1_429 ( .A(_5647_), .B(decoded_rs2_0_bF_buf40_), .C(_5648_), .Y(_5649_) );
MUX2X1 MUX2X1_48 ( .A(_5649_), .B(_5646_), .S(decoded_rs2_1_bF_buf14_), .Y(_5650_) );
AOI21X1 AOI21X1_50 ( .A(_5358__bF_buf2), .B(_5650_), .C(_5348__bF_buf5), .Y(_5651_) );
INVX1 INVX1_318 ( .A(cpuregs_4_[4]), .Y(_5652_) );
NAND2X1 NAND2X1_219 ( .A(cpuregs_5_[4]), .B(decoded_rs2_0_bF_buf39_), .Y(_5653_) );
OAI21X1 OAI21X1_430 ( .A(_5652_), .B(decoded_rs2_0_bF_buf38_), .C(_5653_), .Y(_5654_) );
NAND2X1 NAND2X1_220 ( .A(cpuregs_7_[4]), .B(decoded_rs2_0_bF_buf37_), .Y(_5655_) );
OAI21X1 OAI21X1_431 ( .A(_5278_), .B(decoded_rs2_0_bF_buf36_), .C(_5655_), .Y(_5656_) );
MUX2X1 MUX2X1_49 ( .A(_5656_), .B(_5654_), .S(decoded_rs2_1_bF_buf13_), .Y(_5657_) );
NOR2X1 NOR2X1_251 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_0_[4]), .Y(_5658_) );
OAI21X1 OAI21X1_432 ( .A(_5362__bF_buf12), .B(cpuregs_1_[4]), .C(_5349__bF_buf10), .Y(_5659_) );
NOR2X1 NOR2X1_252 ( .A(_5658_), .B(_5659_), .Y(_5660_) );
INVX1 INVX1_319 ( .A(cpuregs_3_[4]), .Y(_5661_) );
OAI21X1 OAI21X1_433 ( .A(decoded_rs2_0_bF_buf34_), .B(cpuregs_2_[4]), .C(decoded_rs2_1_bF_buf12_), .Y(_5662_) );
AOI21X1 AOI21X1_51 ( .A(decoded_rs2_0_bF_buf33_), .B(_5661_), .C(_5662_), .Y(_5663_) );
OAI21X1 OAI21X1_434 ( .A(_5660_), .B(_5663_), .C(_5358__bF_buf1), .Y(_5664_) );
OAI21X1 OAI21X1_435 ( .A(_5358__bF_buf0), .B(_5657_), .C(_5664_), .Y(_5665_) );
AOI22X1 AOI22X1_11 ( .A(_5643_), .B(_5651_), .C(_5665_), .D(_5348__bF_buf4), .Y(_5666_) );
INVX1 INVX1_320 ( .A(cpuregs_24_[4]), .Y(_5667_) );
OAI21X1 OAI21X1_436 ( .A(_5362__bF_buf11), .B(cpuregs_25_[4]), .C(_5349__bF_buf9), .Y(_5668_) );
AOI21X1 AOI21X1_52 ( .A(_5362__bF_buf10), .B(_5667_), .C(_5668_), .Y(_5669_) );
INVX1 INVX1_321 ( .A(cpuregs_27_[4]), .Y(_5670_) );
OAI21X1 OAI21X1_437 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_26_[4]), .C(decoded_rs2_1_bF_buf11_), .Y(_5671_) );
AOI21X1 AOI21X1_53 ( .A(decoded_rs2_0_bF_buf31_), .B(_5670_), .C(_5671_), .Y(_5672_) );
OAI21X1 OAI21X1_438 ( .A(_5669_), .B(_5672_), .C(_5358__bF_buf12), .Y(_5673_) );
INVX1 INVX1_322 ( .A(cpuregs_28_[4]), .Y(_5674_) );
OAI21X1 OAI21X1_439 ( .A(_5362__bF_buf9), .B(cpuregs_29_[4]), .C(_5349__bF_buf8), .Y(_5675_) );
AOI21X1 AOI21X1_54 ( .A(_5362__bF_buf8), .B(_5674_), .C(_5675_), .Y(_5676_) );
INVX1 INVX1_323 ( .A(cpuregs_31_[4]), .Y(_5677_) );
OAI21X1 OAI21X1_440 ( .A(decoded_rs2_0_bF_buf30_), .B(cpuregs_30_[4]), .C(decoded_rs2_1_bF_buf10_), .Y(_5678_) );
AOI21X1 AOI21X1_55 ( .A(decoded_rs2_0_bF_buf29_), .B(_5677_), .C(_5678_), .Y(_5679_) );
OAI21X1 OAI21X1_441 ( .A(_5676_), .B(_5679_), .C(decoded_rs2_2_bF_buf2_), .Y(_5680_) );
AOI21X1 AOI21X1_56 ( .A(_5673_), .B(_5680_), .C(_5348__bF_buf3), .Y(_5681_) );
INVX1 INVX1_324 ( .A(cpuregs_16_[4]), .Y(_5682_) );
NAND2X1 NAND2X1_221 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_17_[4]), .Y(_5683_) );
OAI21X1 OAI21X1_442 ( .A(_5682_), .B(decoded_rs2_0_bF_buf27_), .C(_5683_), .Y(_5684_) );
INVX1 INVX1_325 ( .A(cpuregs_18_[4]), .Y(_5685_) );
NAND2X1 NAND2X1_222 ( .A(decoded_rs2_0_bF_buf26_), .B(cpuregs_19_[4]), .Y(_5686_) );
OAI21X1 OAI21X1_443 ( .A(_5685_), .B(decoded_rs2_0_bF_buf25_), .C(_5686_), .Y(_5687_) );
MUX2X1 MUX2X1_50 ( .A(_5687_), .B(_5684_), .S(decoded_rs2_1_bF_buf9_), .Y(_5688_) );
INVX1 INVX1_326 ( .A(cpuregs_20_[4]), .Y(_5689_) );
NAND2X1 NAND2X1_223 ( .A(decoded_rs2_0_bF_buf24_), .B(cpuregs_21_[4]), .Y(_5690_) );
OAI21X1 OAI21X1_444 ( .A(_5689_), .B(decoded_rs2_0_bF_buf23_), .C(_5690_), .Y(_5691_) );
INVX1 INVX1_327 ( .A(cpuregs_23_[4]), .Y(_5692_) );
NAND2X1 NAND2X1_224 ( .A(cpuregs_22_[4]), .B(_5362__bF_buf7), .Y(_5693_) );
OAI21X1 OAI21X1_445 ( .A(_5362__bF_buf6), .B(_5692_), .C(_5693_), .Y(_5694_) );
MUX2X1 MUX2X1_51 ( .A(_5694_), .B(_5691_), .S(decoded_rs2_1_bF_buf8_), .Y(_5695_) );
MUX2X1 MUX2X1_52 ( .A(_5695_), .B(_5688_), .S(decoded_rs2_2_bF_buf1_), .Y(_5696_) );
AOI21X1 AOI21X1_57 ( .A(_5348__bF_buf2), .B(_5696_), .C(_5681_), .Y(_5697_) );
NAND2X1 NAND2X1_225 ( .A(decoded_rs2_4_bF_buf2_), .B(_5697_), .Y(_5698_) );
OAI21X1 OAI21X1_446 ( .A(_5384_), .B(_5385_), .C(_5698_), .Y(_5699_) );
AOI21X1 AOI21X1_58 ( .A(_5347_), .B(_5666_), .C(_5699_), .Y(_5700_) );
NOR2X1 NOR2X1_253 ( .A(is_slli_srli_srai), .B(_5700_), .Y(_5701_) );
OAI21X1 OAI21X1_447 ( .A(_4564_), .B(decoded_rs2_4_bF_buf1_), .C(_4575__bF_buf4), .Y(_5702_) );
OAI21X1 OAI21X1_448 ( .A(_5632_), .B(_4577_), .C(_4582_), .Y(_5703_) );
NAND2X1 NAND2X1_226 ( .A(cpu_state_4_), .B(_5703_), .Y(_5704_) );
OAI21X1 OAI21X1_449 ( .A(_5701_), .B(_5702_), .C(_5704_), .Y(_85__4_) );
NOR2X1 NOR2X1_254 ( .A(_4667_), .B(_4632__bF_buf1), .Y(_5705_) );
INVX1 INVX1_328 ( .A(_5705_), .Y(_5706_) );
NOR2X1 NOR2X1_255 ( .A(_4913__bF_buf0), .B(_5706__bF_buf11), .Y(_5707_) );
MUX2X1 MUX2X1_53 ( .A(_4925__bF_buf1), .B(_5368_), .S(_5707__bF_buf3), .Y(_218_) );
MUX2X1 MUX2X1_54 ( .A(_4933__bF_buf1), .B(_5440_), .S(_5707__bF_buf2), .Y(_219_) );
MUX2X1 MUX2X1_55 ( .A(_4940__bF_buf1), .B(_5509_), .S(_5707__bF_buf1), .Y(_220_) );
MUX2X1 MUX2X1_56 ( .A(_4948__bF_buf1), .B(_5581_), .S(_5707__bF_buf0), .Y(_221_) );
MUX2X1 MUX2X1_57 ( .A(_4955__bF_buf1), .B(_5652_), .S(_5707__bF_buf3), .Y(_222_) );
NOR2X1 NOR2X1_256 ( .A(cpuregs_4_[5]), .B(_5707__bF_buf2), .Y(_5708_) );
AOI21X1 AOI21X1_59 ( .A(_4654__bF_buf0), .B(_5707__bF_buf1), .C(_5708_), .Y(_223_) );
INVX1 INVX1_329 ( .A(cpuregs_4_[6]), .Y(_5709_) );
MUX2X1 MUX2X1_58 ( .A(_4664__bF_buf0), .B(_5709_), .S(_5707__bF_buf0), .Y(_224_) );
NOR2X1 NOR2X1_257 ( .A(cpuregs_4_[7]), .B(_5707__bF_buf3), .Y(_5710_) );
AOI21X1 AOI21X1_60 ( .A(_4677__bF_buf0), .B(_5707__bF_buf2), .C(_5710_), .Y(_225_) );
NOR2X1 NOR2X1_258 ( .A(cpuregs_4_[8]), .B(_5707__bF_buf1), .Y(_5711_) );
AOI21X1 AOI21X1_61 ( .A(_5707__bF_buf0), .B(_4685__bF_buf0), .C(_5711_), .Y(_226_) );
NOR2X1 NOR2X1_259 ( .A(cpuregs_4_[9]), .B(_5707__bF_buf3), .Y(_5712_) );
AOI21X1 AOI21X1_62 ( .A(_5707__bF_buf2), .B(_4696__bF_buf0), .C(_5712_), .Y(_227_) );
NOR2X1 NOR2X1_260 ( .A(cpuregs_4_[10]), .B(_5707__bF_buf1), .Y(_5713_) );
AOI21X1 AOI21X1_63 ( .A(_5707__bF_buf0), .B(_4703__bF_buf0), .C(_5713_), .Y(_228_) );
INVX1 INVX1_330 ( .A(cpuregs_4_[11]), .Y(_5714_) );
MUX2X1 MUX2X1_59 ( .A(_4713__bF_buf0), .B(_5714_), .S(_5707__bF_buf3), .Y(_229_) );
INVX1 INVX1_331 ( .A(_5707__bF_buf2), .Y(_5715_) );
OAI21X1 OAI21X1_450 ( .A(_5706__bF_buf10), .B(_4913__bF_buf6), .C(cpuregs_4_[12]), .Y(_5716_) );
OAI21X1 OAI21X1_451 ( .A(_4722__bF_buf0), .B(_5715__bF_buf3), .C(_5716_), .Y(_230_) );
OAI21X1 OAI21X1_452 ( .A(_5706__bF_buf9), .B(_4913__bF_buf5), .C(cpuregs_4_[13]), .Y(_5717_) );
OAI21X1 OAI21X1_453 ( .A(_4731__bF_buf0), .B(_5715__bF_buf2), .C(_5717_), .Y(_231_) );
OAI21X1 OAI21X1_454 ( .A(_5706__bF_buf8), .B(_4913__bF_buf4), .C(cpuregs_4_[14]), .Y(_5718_) );
OAI21X1 OAI21X1_455 ( .A(_4740__bF_buf0), .B(_5715__bF_buf1), .C(_5718_), .Y(_232_) );
OAI21X1 OAI21X1_456 ( .A(_5706__bF_buf7), .B(_4913__bF_buf3), .C(cpuregs_4_[15]), .Y(_5719_) );
OAI21X1 OAI21X1_457 ( .A(_4747__bF_buf0), .B(_5715__bF_buf0), .C(_5719_), .Y(_233_) );
OAI21X1 OAI21X1_458 ( .A(_5706__bF_buf6), .B(_4913__bF_buf2), .C(cpuregs_4_[16]), .Y(_5720_) );
OAI21X1 OAI21X1_459 ( .A(_4755__bF_buf0), .B(_5715__bF_buf3), .C(_5720_), .Y(_234_) );
OAI21X1 OAI21X1_460 ( .A(_5706__bF_buf5), .B(_4913__bF_buf1), .C(cpuregs_4_[17]), .Y(_5721_) );
OAI21X1 OAI21X1_461 ( .A(_4763__bF_buf0), .B(_5715__bF_buf2), .C(_5721_), .Y(_235_) );
OAI21X1 OAI21X1_462 ( .A(_5706__bF_buf4), .B(_4913__bF_buf0), .C(cpuregs_4_[18]), .Y(_5722_) );
OAI21X1 OAI21X1_463 ( .A(_4783__bF_buf0), .B(_5715__bF_buf1), .C(_5722_), .Y(_236_) );
OAI21X1 OAI21X1_464 ( .A(_5706__bF_buf3), .B(_4913__bF_buf6), .C(cpuregs_4_[19]), .Y(_5723_) );
OAI21X1 OAI21X1_465 ( .A(_4793__bF_buf0), .B(_5715__bF_buf0), .C(_5723_), .Y(_237_) );
OAI21X1 OAI21X1_466 ( .A(_5706__bF_buf2), .B(_4913__bF_buf5), .C(cpuregs_4_[20]), .Y(_5724_) );
OAI21X1 OAI21X1_467 ( .A(_4806__bF_buf0), .B(_5715__bF_buf3), .C(_5724_), .Y(_238_) );
OAI21X1 OAI21X1_468 ( .A(_5706__bF_buf1), .B(_4913__bF_buf4), .C(cpuregs_4_[21]), .Y(_5725_) );
OAI21X1 OAI21X1_469 ( .A(_4816__bF_buf0), .B(_5715__bF_buf2), .C(_5725_), .Y(_239_) );
OAI21X1 OAI21X1_470 ( .A(_5706__bF_buf0), .B(_4913__bF_buf3), .C(cpuregs_4_[22]), .Y(_5726_) );
OAI21X1 OAI21X1_471 ( .A(_4824__bF_buf0), .B(_5715__bF_buf1), .C(_5726_), .Y(_240_) );
OAI21X1 OAI21X1_472 ( .A(_5706__bF_buf11), .B(_4913__bF_buf2), .C(cpuregs_4_[23]), .Y(_5727_) );
OAI21X1 OAI21X1_473 ( .A(_4833__bF_buf0), .B(_5715__bF_buf0), .C(_5727_), .Y(_241_) );
OAI21X1 OAI21X1_474 ( .A(_5706__bF_buf10), .B(_4913__bF_buf1), .C(cpuregs_4_[24]), .Y(_5728_) );
OAI21X1 OAI21X1_475 ( .A(_4845__bF_buf0), .B(_5715__bF_buf3), .C(_5728_), .Y(_242_) );
OAI21X1 OAI21X1_476 ( .A(_5706__bF_buf9), .B(_4913__bF_buf0), .C(cpuregs_4_[25]), .Y(_5729_) );
OAI21X1 OAI21X1_477 ( .A(_4854__bF_buf0), .B(_5715__bF_buf2), .C(_5729_), .Y(_243_) );
OAI21X1 OAI21X1_478 ( .A(_5706__bF_buf8), .B(_4913__bF_buf6), .C(cpuregs_4_[26]), .Y(_5730_) );
OAI21X1 OAI21X1_479 ( .A(_4863__bF_buf0), .B(_5715__bF_buf1), .C(_5730_), .Y(_244_) );
OAI21X1 OAI21X1_480 ( .A(_5706__bF_buf7), .B(_4913__bF_buf5), .C(cpuregs_4_[27]), .Y(_5731_) );
OAI21X1 OAI21X1_481 ( .A(_4871__bF_buf0), .B(_5715__bF_buf0), .C(_5731_), .Y(_245_) );
OAI21X1 OAI21X1_482 ( .A(_5706__bF_buf6), .B(_4913__bF_buf4), .C(cpuregs_4_[28]), .Y(_5732_) );
OAI21X1 OAI21X1_483 ( .A(_4884__bF_buf0), .B(_5715__bF_buf3), .C(_5732_), .Y(_246_) );
OAI21X1 OAI21X1_484 ( .A(_5706__bF_buf5), .B(_4913__bF_buf3), .C(cpuregs_4_[29]), .Y(_5733_) );
OAI21X1 OAI21X1_485 ( .A(_4893__bF_buf0), .B(_5715__bF_buf2), .C(_5733_), .Y(_247_) );
OAI21X1 OAI21X1_486 ( .A(_5706__bF_buf4), .B(_4913__bF_buf2), .C(cpuregs_4_[30]), .Y(_5734_) );
OAI21X1 OAI21X1_487 ( .A(_4901__bF_buf0), .B(_5715__bF_buf1), .C(_5734_), .Y(_248_) );
OAI21X1 OAI21X1_488 ( .A(_5706__bF_buf3), .B(_4913__bF_buf1), .C(cpuregs_4_[31]), .Y(_5735_) );
OAI21X1 OAI21X1_489 ( .A(_4910__bF_buf0), .B(_5715__bF_buf0), .C(_5735_), .Y(_249_) );
INVX1 INVX1_332 ( .A(decoded_rd_0_), .Y(_5736_) );
NOR2X1 NOR2X1_261 ( .A(is_beq_bne_blt_bge_bltu_bgeu), .B(_4555_), .Y(_5737_) );
OAI21X1 OAI21X1_490 ( .A(cpu_state_3_bF_buf4_), .B(cpu_state_1_bF_buf2_), .C(resetn_bF_buf4), .Y(_5738_) );
NOR2X1 NOR2X1_262 ( .A(_5738_), .B(_5737_), .Y(_5739_) );
OAI22X1 OAI22X1_7 ( .A(_5736_), .B(_4475_), .C(_5739_), .D(_4915_), .Y(_67__0_) );
INVX1 INVX1_333 ( .A(decoded_rd_1_), .Y(_5740_) );
OAI22X1 OAI22X1_8 ( .A(_5740_), .B(_4475_), .C(_5739_), .D(_4914_), .Y(_67__1_) );
INVX1 INVX1_334 ( .A(decoded_rd_2_), .Y(_5741_) );
OAI22X1 OAI22X1_9 ( .A(_5741_), .B(_4475_), .C(_5739_), .D(_4911_), .Y(_67__2_) );
INVX1 INVX1_335 ( .A(decoded_rd_3_), .Y(_5742_) );
OAI22X1 OAI22X1_10 ( .A(_5742_), .B(_4475_), .C(_5739_), .D(_4633_), .Y(_67__3_) );
INVX1 INVX1_336 ( .A(latched_rd_4_), .Y(_5743_) );
INVX1 INVX1_337 ( .A(decoded_rd_4_), .Y(_5744_) );
OAI22X1 OAI22X1_11 ( .A(_5744_), .B(_4475_), .C(_5739_), .D(_5743_), .Y(_67__4_) );
INVX1 INVX1_338 ( .A(_4917__bF_buf10), .Y(_5745_) );
NAND2X1 NAND2X1_227 ( .A(_4627_), .B(_5745_), .Y(_5746_) );
NAND2X1 NAND2X1_228 ( .A(cpuregs_3_[0]), .B(_5746__bF_buf7), .Y(_5747_) );
OAI21X1 OAI21X1_491 ( .A(_4925__bF_buf0), .B(_5746__bF_buf6), .C(_5747_), .Y(_250_) );
NAND2X1 NAND2X1_229 ( .A(cpuregs_3_[1]), .B(_5746__bF_buf5), .Y(_5748_) );
OAI21X1 OAI21X1_492 ( .A(_4933__bF_buf0), .B(_5746__bF_buf4), .C(_5748_), .Y(_251_) );
NAND2X1 NAND2X1_230 ( .A(cpuregs_3_[2]), .B(_5746__bF_buf3), .Y(_5749_) );
OAI21X1 OAI21X1_493 ( .A(_4940__bF_buf0), .B(_5746__bF_buf2), .C(_5749_), .Y(_252_) );
NAND2X1 NAND2X1_231 ( .A(cpuregs_3_[3]), .B(_5746__bF_buf1), .Y(_5750_) );
OAI21X1 OAI21X1_494 ( .A(_4948__bF_buf0), .B(_5746__bF_buf0), .C(_5750_), .Y(_253_) );
NAND2X1 NAND2X1_232 ( .A(cpuregs_3_[4]), .B(_5746__bF_buf7), .Y(_5751_) );
OAI21X1 OAI21X1_495 ( .A(_4955__bF_buf0), .B(_5746__bF_buf6), .C(_5751_), .Y(_254_) );
NAND2X1 NAND2X1_233 ( .A(cpuregs_3_[5]), .B(_5746__bF_buf5), .Y(_5752_) );
OAI21X1 OAI21X1_496 ( .A(_4654__bF_buf4), .B(_5746__bF_buf4), .C(_5752_), .Y(_255_) );
NAND2X1 NAND2X1_234 ( .A(cpuregs_3_[6]), .B(_5746__bF_buf3), .Y(_5753_) );
OAI21X1 OAI21X1_497 ( .A(_4664__bF_buf4), .B(_5746__bF_buf2), .C(_5753_), .Y(_256_) );
NAND2X1 NAND2X1_235 ( .A(cpuregs_3_[7]), .B(_5746__bF_buf1), .Y(_5754_) );
OAI21X1 OAI21X1_498 ( .A(_4677__bF_buf4), .B(_5746__bF_buf0), .C(_5754_), .Y(_257_) );
NAND2X1 NAND2X1_236 ( .A(cpuregs_3_[8]), .B(_5746__bF_buf7), .Y(_5755_) );
OAI21X1 OAI21X1_499 ( .A(_4685__bF_buf4), .B(_5746__bF_buf6), .C(_5755_), .Y(_258_) );
NAND2X1 NAND2X1_237 ( .A(cpuregs_3_[9]), .B(_5746__bF_buf5), .Y(_5756_) );
OAI21X1 OAI21X1_500 ( .A(_4696__bF_buf4), .B(_5746__bF_buf4), .C(_5756_), .Y(_259_) );
NAND2X1 NAND2X1_238 ( .A(cpuregs_3_[10]), .B(_5746__bF_buf3), .Y(_5757_) );
OAI21X1 OAI21X1_501 ( .A(_4703__bF_buf4), .B(_5746__bF_buf2), .C(_5757_), .Y(_260_) );
NAND2X1 NAND2X1_239 ( .A(cpuregs_3_[11]), .B(_5746__bF_buf1), .Y(_5758_) );
OAI21X1 OAI21X1_502 ( .A(_4713__bF_buf4), .B(_5746__bF_buf0), .C(_5758_), .Y(_261_) );
NAND2X1 NAND2X1_240 ( .A(cpuregs_3_[12]), .B(_5746__bF_buf7), .Y(_5759_) );
OAI21X1 OAI21X1_503 ( .A(_4722__bF_buf4), .B(_5746__bF_buf6), .C(_5759_), .Y(_262_) );
NAND2X1 NAND2X1_241 ( .A(cpuregs_3_[13]), .B(_5746__bF_buf5), .Y(_5760_) );
OAI21X1 OAI21X1_504 ( .A(_4731__bF_buf4), .B(_5746__bF_buf4), .C(_5760_), .Y(_263_) );
NAND2X1 NAND2X1_242 ( .A(cpuregs_3_[14]), .B(_5746__bF_buf3), .Y(_5761_) );
OAI21X1 OAI21X1_505 ( .A(_4740__bF_buf4), .B(_5746__bF_buf2), .C(_5761_), .Y(_264_) );
NAND2X1 NAND2X1_243 ( .A(cpuregs_3_[15]), .B(_5746__bF_buf1), .Y(_5762_) );
OAI21X1 OAI21X1_506 ( .A(_4747__bF_buf4), .B(_5746__bF_buf0), .C(_5762_), .Y(_265_) );
NAND2X1 NAND2X1_244 ( .A(cpuregs_3_[16]), .B(_5746__bF_buf7), .Y(_5763_) );
OAI21X1 OAI21X1_507 ( .A(_4755__bF_buf4), .B(_5746__bF_buf6), .C(_5763_), .Y(_266_) );
NAND2X1 NAND2X1_245 ( .A(cpuregs_3_[17]), .B(_5746__bF_buf5), .Y(_5764_) );
OAI21X1 OAI21X1_508 ( .A(_4763__bF_buf4), .B(_5746__bF_buf4), .C(_5764_), .Y(_267_) );
NAND2X1 NAND2X1_246 ( .A(cpuregs_3_[18]), .B(_5746__bF_buf3), .Y(_5765_) );
OAI21X1 OAI21X1_509 ( .A(_4783__bF_buf4), .B(_5746__bF_buf2), .C(_5765_), .Y(_268_) );
NAND2X1 NAND2X1_247 ( .A(cpuregs_3_[19]), .B(_5746__bF_buf1), .Y(_5766_) );
OAI21X1 OAI21X1_510 ( .A(_4793__bF_buf4), .B(_5746__bF_buf0), .C(_5766_), .Y(_269_) );
NAND2X1 NAND2X1_248 ( .A(cpuregs_3_[20]), .B(_5746__bF_buf7), .Y(_5767_) );
OAI21X1 OAI21X1_511 ( .A(_4806__bF_buf4), .B(_5746__bF_buf6), .C(_5767_), .Y(_270_) );
NAND2X1 NAND2X1_249 ( .A(cpuregs_3_[21]), .B(_5746__bF_buf5), .Y(_5768_) );
OAI21X1 OAI21X1_512 ( .A(_4816__bF_buf4), .B(_5746__bF_buf4), .C(_5768_), .Y(_271_) );
NAND2X1 NAND2X1_250 ( .A(cpuregs_3_[22]), .B(_5746__bF_buf3), .Y(_5769_) );
OAI21X1 OAI21X1_513 ( .A(_4824__bF_buf4), .B(_5746__bF_buf2), .C(_5769_), .Y(_272_) );
NAND2X1 NAND2X1_251 ( .A(cpuregs_3_[23]), .B(_5746__bF_buf1), .Y(_5770_) );
OAI21X1 OAI21X1_514 ( .A(_4833__bF_buf4), .B(_5746__bF_buf0), .C(_5770_), .Y(_273_) );
NAND2X1 NAND2X1_252 ( .A(cpuregs_3_[24]), .B(_5746__bF_buf7), .Y(_5771_) );
OAI21X1 OAI21X1_515 ( .A(_4845__bF_buf4), .B(_5746__bF_buf6), .C(_5771_), .Y(_274_) );
NAND2X1 NAND2X1_253 ( .A(cpuregs_3_[25]), .B(_5746__bF_buf5), .Y(_5772_) );
OAI21X1 OAI21X1_516 ( .A(_4854__bF_buf4), .B(_5746__bF_buf4), .C(_5772_), .Y(_275_) );
NAND2X1 NAND2X1_254 ( .A(cpuregs_3_[26]), .B(_5746__bF_buf3), .Y(_5773_) );
OAI21X1 OAI21X1_517 ( .A(_4863__bF_buf4), .B(_5746__bF_buf2), .C(_5773_), .Y(_276_) );
NAND2X1 NAND2X1_255 ( .A(cpuregs_3_[27]), .B(_5746__bF_buf1), .Y(_5774_) );
OAI21X1 OAI21X1_518 ( .A(_4871__bF_buf4), .B(_5746__bF_buf0), .C(_5774_), .Y(_277_) );
NAND2X1 NAND2X1_256 ( .A(cpuregs_3_[28]), .B(_5746__bF_buf7), .Y(_5775_) );
OAI21X1 OAI21X1_519 ( .A(_4884__bF_buf4), .B(_5746__bF_buf6), .C(_5775_), .Y(_278_) );
NAND2X1 NAND2X1_257 ( .A(cpuregs_3_[29]), .B(_5746__bF_buf5), .Y(_5776_) );
OAI21X1 OAI21X1_520 ( .A(_4893__bF_buf4), .B(_5746__bF_buf4), .C(_5776_), .Y(_279_) );
NAND2X1 NAND2X1_258 ( .A(cpuregs_3_[30]), .B(_5746__bF_buf3), .Y(_5777_) );
OAI21X1 OAI21X1_521 ( .A(_4901__bF_buf4), .B(_5746__bF_buf2), .C(_5777_), .Y(_280_) );
NAND2X1 NAND2X1_259 ( .A(cpuregs_3_[31]), .B(_5746__bF_buf1), .Y(_5778_) );
OAI21X1 OAI21X1_522 ( .A(_4910__bF_buf4), .B(_5746__bF_buf0), .C(_5778_), .Y(_281_) );
INVX1 INVX1_339 ( .A(_5281__bF_buf9), .Y(_5779_) );
NAND2X1 NAND2X1_260 ( .A(_4627_), .B(_5779_), .Y(_5780_) );
NAND2X1 NAND2X1_261 ( .A(cpuregs_2_[0]), .B(_5780__bF_buf7), .Y(_5781_) );
OAI21X1 OAI21X1_523 ( .A(_4925__bF_buf4), .B(_5780__bF_buf6), .C(_5781_), .Y(_282_) );
NAND2X1 NAND2X1_262 ( .A(cpuregs_2_[1]), .B(_5780__bF_buf5), .Y(_5782_) );
OAI21X1 OAI21X1_524 ( .A(_4933__bF_buf4), .B(_5780__bF_buf4), .C(_5782_), .Y(_283_) );
NAND2X1 NAND2X1_263 ( .A(cpuregs_2_[2]), .B(_5780__bF_buf3), .Y(_5783_) );
OAI21X1 OAI21X1_525 ( .A(_4940__bF_buf4), .B(_5780__bF_buf2), .C(_5783_), .Y(_284_) );
NAND2X1 NAND2X1_264 ( .A(cpuregs_2_[3]), .B(_5780__bF_buf1), .Y(_5784_) );
OAI21X1 OAI21X1_526 ( .A(_4948__bF_buf4), .B(_5780__bF_buf0), .C(_5784_), .Y(_285_) );
NAND2X1 NAND2X1_265 ( .A(cpuregs_2_[4]), .B(_5780__bF_buf7), .Y(_5785_) );
OAI21X1 OAI21X1_527 ( .A(_4955__bF_buf4), .B(_5780__bF_buf6), .C(_5785_), .Y(_286_) );
NAND2X1 NAND2X1_266 ( .A(cpuregs_2_[5]), .B(_5780__bF_buf5), .Y(_5786_) );
OAI21X1 OAI21X1_528 ( .A(_4654__bF_buf3), .B(_5780__bF_buf4), .C(_5786_), .Y(_287_) );
NAND2X1 NAND2X1_267 ( .A(cpuregs_2_[6]), .B(_5780__bF_buf3), .Y(_5787_) );
OAI21X1 OAI21X1_529 ( .A(_4664__bF_buf3), .B(_5780__bF_buf2), .C(_5787_), .Y(_288_) );
NAND2X1 NAND2X1_268 ( .A(cpuregs_2_[7]), .B(_5780__bF_buf1), .Y(_5788_) );
OAI21X1 OAI21X1_530 ( .A(_4677__bF_buf3), .B(_5780__bF_buf0), .C(_5788_), .Y(_289_) );
NAND2X1 NAND2X1_269 ( .A(cpuregs_2_[8]), .B(_5780__bF_buf7), .Y(_5789_) );
OAI21X1 OAI21X1_531 ( .A(_4685__bF_buf3), .B(_5780__bF_buf6), .C(_5789_), .Y(_290_) );
NAND2X1 NAND2X1_270 ( .A(cpuregs_2_[9]), .B(_5780__bF_buf5), .Y(_5790_) );
OAI21X1 OAI21X1_532 ( .A(_4696__bF_buf3), .B(_5780__bF_buf4), .C(_5790_), .Y(_291_) );
NAND2X1 NAND2X1_271 ( .A(cpuregs_2_[10]), .B(_5780__bF_buf3), .Y(_5791_) );
OAI21X1 OAI21X1_533 ( .A(_4703__bF_buf3), .B(_5780__bF_buf2), .C(_5791_), .Y(_292_) );
NAND2X1 NAND2X1_272 ( .A(cpuregs_2_[11]), .B(_5780__bF_buf1), .Y(_5792_) );
OAI21X1 OAI21X1_534 ( .A(_4713__bF_buf3), .B(_5780__bF_buf0), .C(_5792_), .Y(_293_) );
NAND2X1 NAND2X1_273 ( .A(cpuregs_2_[12]), .B(_5780__bF_buf7), .Y(_5793_) );
OAI21X1 OAI21X1_535 ( .A(_4722__bF_buf3), .B(_5780__bF_buf6), .C(_5793_), .Y(_294_) );
NAND2X1 NAND2X1_274 ( .A(cpuregs_2_[13]), .B(_5780__bF_buf5), .Y(_5794_) );
OAI21X1 OAI21X1_536 ( .A(_4731__bF_buf3), .B(_5780__bF_buf4), .C(_5794_), .Y(_295_) );
NAND2X1 NAND2X1_275 ( .A(cpuregs_2_[14]), .B(_5780__bF_buf3), .Y(_5795_) );
OAI21X1 OAI21X1_537 ( .A(_4740__bF_buf3), .B(_5780__bF_buf2), .C(_5795_), .Y(_296_) );
NAND2X1 NAND2X1_276 ( .A(cpuregs_2_[15]), .B(_5780__bF_buf1), .Y(_5796_) );
OAI21X1 OAI21X1_538 ( .A(_4747__bF_buf3), .B(_5780__bF_buf0), .C(_5796_), .Y(_297_) );
NAND2X1 NAND2X1_277 ( .A(cpuregs_2_[16]), .B(_5780__bF_buf7), .Y(_5797_) );
OAI21X1 OAI21X1_539 ( .A(_4755__bF_buf3), .B(_5780__bF_buf6), .C(_5797_), .Y(_298_) );
NAND2X1 NAND2X1_278 ( .A(cpuregs_2_[17]), .B(_5780__bF_buf5), .Y(_5798_) );
OAI21X1 OAI21X1_540 ( .A(_4763__bF_buf3), .B(_5780__bF_buf4), .C(_5798_), .Y(_299_) );
NAND2X1 NAND2X1_279 ( .A(cpuregs_2_[18]), .B(_5780__bF_buf3), .Y(_5799_) );
OAI21X1 OAI21X1_541 ( .A(_4783__bF_buf3), .B(_5780__bF_buf2), .C(_5799_), .Y(_300_) );
NAND2X1 NAND2X1_280 ( .A(cpuregs_2_[19]), .B(_5780__bF_buf1), .Y(_5800_) );
OAI21X1 OAI21X1_542 ( .A(_4793__bF_buf3), .B(_5780__bF_buf0), .C(_5800_), .Y(_301_) );
NAND2X1 NAND2X1_281 ( .A(cpuregs_2_[20]), .B(_5780__bF_buf7), .Y(_5801_) );
OAI21X1 OAI21X1_543 ( .A(_4806__bF_buf3), .B(_5780__bF_buf6), .C(_5801_), .Y(_302_) );
NAND2X1 NAND2X1_282 ( .A(cpuregs_2_[21]), .B(_5780__bF_buf5), .Y(_5802_) );
OAI21X1 OAI21X1_544 ( .A(_4816__bF_buf3), .B(_5780__bF_buf4), .C(_5802_), .Y(_303_) );
NAND2X1 NAND2X1_283 ( .A(cpuregs_2_[22]), .B(_5780__bF_buf3), .Y(_5803_) );
OAI21X1 OAI21X1_545 ( .A(_4824__bF_buf3), .B(_5780__bF_buf2), .C(_5803_), .Y(_304_) );
NAND2X1 NAND2X1_284 ( .A(cpuregs_2_[23]), .B(_5780__bF_buf1), .Y(_5804_) );
OAI21X1 OAI21X1_546 ( .A(_4833__bF_buf3), .B(_5780__bF_buf0), .C(_5804_), .Y(_305_) );
NAND2X1 NAND2X1_285 ( .A(cpuregs_2_[24]), .B(_5780__bF_buf7), .Y(_5805_) );
OAI21X1 OAI21X1_547 ( .A(_4845__bF_buf3), .B(_5780__bF_buf6), .C(_5805_), .Y(_306_) );
NAND2X1 NAND2X1_286 ( .A(cpuregs_2_[25]), .B(_5780__bF_buf5), .Y(_5806_) );
OAI21X1 OAI21X1_548 ( .A(_4854__bF_buf3), .B(_5780__bF_buf4), .C(_5806_), .Y(_307_) );
NAND2X1 NAND2X1_287 ( .A(cpuregs_2_[26]), .B(_5780__bF_buf3), .Y(_5807_) );
OAI21X1 OAI21X1_549 ( .A(_4863__bF_buf3), .B(_5780__bF_buf2), .C(_5807_), .Y(_308_) );
NAND2X1 NAND2X1_288 ( .A(cpuregs_2_[27]), .B(_5780__bF_buf1), .Y(_5808_) );
OAI21X1 OAI21X1_550 ( .A(_4871__bF_buf3), .B(_5780__bF_buf0), .C(_5808_), .Y(_309_) );
NAND2X1 NAND2X1_289 ( .A(cpuregs_2_[28]), .B(_5780__bF_buf7), .Y(_5809_) );
OAI21X1 OAI21X1_551 ( .A(_4884__bF_buf3), .B(_5780__bF_buf6), .C(_5809_), .Y(_310_) );
NAND2X1 NAND2X1_290 ( .A(cpuregs_2_[29]), .B(_5780__bF_buf5), .Y(_5810_) );
OAI21X1 OAI21X1_552 ( .A(_4893__bF_buf3), .B(_5780__bF_buf4), .C(_5810_), .Y(_311_) );
NAND2X1 NAND2X1_291 ( .A(cpuregs_2_[30]), .B(_5780__bF_buf3), .Y(_5811_) );
OAI21X1 OAI21X1_553 ( .A(_4901__bF_buf3), .B(_5780__bF_buf2), .C(_5811_), .Y(_312_) );
NAND2X1 NAND2X1_292 ( .A(cpuregs_2_[31]), .B(_5780__bF_buf1), .Y(_5812_) );
OAI21X1 OAI21X1_554 ( .A(_4910__bF_buf3), .B(_5780__bF_buf0), .C(_5812_), .Y(_313_) );
AND2X2 AND2X2_22 ( .A(_4475_), .B(latched_compr), .Y(_64_) );
NAND2X1 NAND2X1_293 ( .A(_4627_), .B(_5313_), .Y(_5813_) );
NAND2X1 NAND2X1_294 ( .A(cpuregs_1_[0]), .B(_5813__bF_buf7), .Y(_5814_) );
OAI21X1 OAI21X1_555 ( .A(_4925__bF_buf3), .B(_5813__bF_buf6), .C(_5814_), .Y(_314_) );
NAND2X1 NAND2X1_295 ( .A(cpuregs_1_[1]), .B(_5813__bF_buf5), .Y(_5815_) );
OAI21X1 OAI21X1_556 ( .A(_4933__bF_buf3), .B(_5813__bF_buf4), .C(_5815_), .Y(_315_) );
NAND2X1 NAND2X1_296 ( .A(cpuregs_1_[2]), .B(_5813__bF_buf3), .Y(_5816_) );
OAI21X1 OAI21X1_557 ( .A(_4940__bF_buf3), .B(_5813__bF_buf2), .C(_5816_), .Y(_316_) );
NAND2X1 NAND2X1_297 ( .A(cpuregs_1_[3]), .B(_5813__bF_buf1), .Y(_5817_) );
OAI21X1 OAI21X1_558 ( .A(_4948__bF_buf3), .B(_5813__bF_buf0), .C(_5817_), .Y(_317_) );
NAND2X1 NAND2X1_298 ( .A(cpuregs_1_[4]), .B(_5813__bF_buf7), .Y(_5818_) );
OAI21X1 OAI21X1_559 ( .A(_4955__bF_buf3), .B(_5813__bF_buf6), .C(_5818_), .Y(_318_) );
NAND2X1 NAND2X1_299 ( .A(cpuregs_1_[5]), .B(_5813__bF_buf5), .Y(_5819_) );
OAI21X1 OAI21X1_560 ( .A(_4654__bF_buf2), .B(_5813__bF_buf4), .C(_5819_), .Y(_319_) );
NAND2X1 NAND2X1_300 ( .A(cpuregs_1_[6]), .B(_5813__bF_buf3), .Y(_5820_) );
OAI21X1 OAI21X1_561 ( .A(_4664__bF_buf2), .B(_5813__bF_buf2), .C(_5820_), .Y(_320_) );
NAND2X1 NAND2X1_301 ( .A(cpuregs_1_[7]), .B(_5813__bF_buf1), .Y(_5821_) );
OAI21X1 OAI21X1_562 ( .A(_4677__bF_buf2), .B(_5813__bF_buf0), .C(_5821_), .Y(_321_) );
NAND2X1 NAND2X1_302 ( .A(cpuregs_1_[8]), .B(_5813__bF_buf7), .Y(_5822_) );
OAI21X1 OAI21X1_563 ( .A(_4685__bF_buf2), .B(_5813__bF_buf6), .C(_5822_), .Y(_322_) );
NAND2X1 NAND2X1_303 ( .A(cpuregs_1_[9]), .B(_5813__bF_buf5), .Y(_5823_) );
OAI21X1 OAI21X1_564 ( .A(_4696__bF_buf2), .B(_5813__bF_buf4), .C(_5823_), .Y(_323_) );
NAND2X1 NAND2X1_304 ( .A(cpuregs_1_[10]), .B(_5813__bF_buf3), .Y(_5824_) );
OAI21X1 OAI21X1_565 ( .A(_4703__bF_buf2), .B(_5813__bF_buf2), .C(_5824_), .Y(_324_) );
NAND2X1 NAND2X1_305 ( .A(cpuregs_1_[11]), .B(_5813__bF_buf1), .Y(_5825_) );
OAI21X1 OAI21X1_566 ( .A(_4713__bF_buf2), .B(_5813__bF_buf0), .C(_5825_), .Y(_325_) );
NAND2X1 NAND2X1_306 ( .A(cpuregs_1_[12]), .B(_5813__bF_buf7), .Y(_5826_) );
OAI21X1 OAI21X1_567 ( .A(_4722__bF_buf2), .B(_5813__bF_buf6), .C(_5826_), .Y(_326_) );
NAND2X1 NAND2X1_307 ( .A(cpuregs_1_[13]), .B(_5813__bF_buf5), .Y(_5827_) );
OAI21X1 OAI21X1_568 ( .A(_4731__bF_buf2), .B(_5813__bF_buf4), .C(_5827_), .Y(_327_) );
NAND2X1 NAND2X1_308 ( .A(cpuregs_1_[14]), .B(_5813__bF_buf3), .Y(_5828_) );
OAI21X1 OAI21X1_569 ( .A(_4740__bF_buf2), .B(_5813__bF_buf2), .C(_5828_), .Y(_328_) );
NAND2X1 NAND2X1_309 ( .A(cpuregs_1_[15]), .B(_5813__bF_buf1), .Y(_5829_) );
OAI21X1 OAI21X1_570 ( .A(_4747__bF_buf2), .B(_5813__bF_buf0), .C(_5829_), .Y(_329_) );
NAND2X1 NAND2X1_310 ( .A(cpuregs_1_[16]), .B(_5813__bF_buf7), .Y(_5830_) );
OAI21X1 OAI21X1_571 ( .A(_4755__bF_buf2), .B(_5813__bF_buf6), .C(_5830_), .Y(_330_) );
NAND2X1 NAND2X1_311 ( .A(cpuregs_1_[17]), .B(_5813__bF_buf5), .Y(_5831_) );
OAI21X1 OAI21X1_572 ( .A(_4763__bF_buf2), .B(_5813__bF_buf4), .C(_5831_), .Y(_331_) );
NAND2X1 NAND2X1_312 ( .A(cpuregs_1_[18]), .B(_5813__bF_buf3), .Y(_5832_) );
OAI21X1 OAI21X1_573 ( .A(_4783__bF_buf2), .B(_5813__bF_buf2), .C(_5832_), .Y(_332_) );
NAND2X1 NAND2X1_313 ( .A(cpuregs_1_[19]), .B(_5813__bF_buf1), .Y(_5833_) );
OAI21X1 OAI21X1_574 ( .A(_4793__bF_buf2), .B(_5813__bF_buf0), .C(_5833_), .Y(_333_) );
NAND2X1 NAND2X1_314 ( .A(cpuregs_1_[20]), .B(_5813__bF_buf7), .Y(_5834_) );
OAI21X1 OAI21X1_575 ( .A(_4806__bF_buf2), .B(_5813__bF_buf6), .C(_5834_), .Y(_334_) );
NAND2X1 NAND2X1_315 ( .A(cpuregs_1_[21]), .B(_5813__bF_buf5), .Y(_5835_) );
OAI21X1 OAI21X1_576 ( .A(_4816__bF_buf2), .B(_5813__bF_buf4), .C(_5835_), .Y(_335_) );
NAND2X1 NAND2X1_316 ( .A(cpuregs_1_[22]), .B(_5813__bF_buf3), .Y(_5836_) );
OAI21X1 OAI21X1_577 ( .A(_4824__bF_buf2), .B(_5813__bF_buf2), .C(_5836_), .Y(_336_) );
NAND2X1 NAND2X1_317 ( .A(cpuregs_1_[23]), .B(_5813__bF_buf1), .Y(_5837_) );
OAI21X1 OAI21X1_578 ( .A(_4833__bF_buf2), .B(_5813__bF_buf0), .C(_5837_), .Y(_337_) );
NAND2X1 NAND2X1_318 ( .A(cpuregs_1_[24]), .B(_5813__bF_buf7), .Y(_5838_) );
OAI21X1 OAI21X1_579 ( .A(_4845__bF_buf2), .B(_5813__bF_buf6), .C(_5838_), .Y(_338_) );
NAND2X1 NAND2X1_319 ( .A(cpuregs_1_[25]), .B(_5813__bF_buf5), .Y(_5839_) );
OAI21X1 OAI21X1_580 ( .A(_4854__bF_buf2), .B(_5813__bF_buf4), .C(_5839_), .Y(_339_) );
NAND2X1 NAND2X1_320 ( .A(cpuregs_1_[26]), .B(_5813__bF_buf3), .Y(_5840_) );
OAI21X1 OAI21X1_581 ( .A(_4863__bF_buf2), .B(_5813__bF_buf2), .C(_5840_), .Y(_340_) );
NAND2X1 NAND2X1_321 ( .A(cpuregs_1_[27]), .B(_5813__bF_buf1), .Y(_5841_) );
OAI21X1 OAI21X1_582 ( .A(_4871__bF_buf2), .B(_5813__bF_buf0), .C(_5841_), .Y(_341_) );
NAND2X1 NAND2X1_322 ( .A(cpuregs_1_[28]), .B(_5813__bF_buf7), .Y(_5842_) );
OAI21X1 OAI21X1_583 ( .A(_4884__bF_buf2), .B(_5813__bF_buf6), .C(_5842_), .Y(_342_) );
NAND2X1 NAND2X1_323 ( .A(cpuregs_1_[29]), .B(_5813__bF_buf5), .Y(_5843_) );
OAI21X1 OAI21X1_584 ( .A(_4893__bF_buf2), .B(_5813__bF_buf4), .C(_5843_), .Y(_343_) );
NAND2X1 NAND2X1_324 ( .A(cpuregs_1_[30]), .B(_5813__bF_buf3), .Y(_5844_) );
OAI21X1 OAI21X1_585 ( .A(_4901__bF_buf2), .B(_5813__bF_buf2), .C(_5844_), .Y(_344_) );
NAND2X1 NAND2X1_325 ( .A(cpuregs_1_[31]), .B(_5813__bF_buf1), .Y(_5845_) );
OAI21X1 OAI21X1_586 ( .A(_4910__bF_buf2), .B(_5813__bF_buf0), .C(_5845_), .Y(_345_) );
OAI21X1 OAI21X1_587 ( .A(_4475_), .B(_4611_), .C(mem_do_prefetch_bF_buf0), .Y(_5846_) );
INVX1 INVX1_340 ( .A(instr_jalr), .Y(_5847_) );
NAND2X1 NAND2X1_326 ( .A(_5847_), .B(_4612_), .Y(_5848_) );
AOI21X1 AOI21X1_64 ( .A(_5846_), .B(_5848_), .C(_4455_), .Y(_71_) );
INVX1 INVX1_341 ( .A(_4552_), .Y(_5849_) );
NOR2X1 NOR2X1_263 ( .A(_5849__bF_buf4), .B(_5419_), .Y(_5850_) );
OAI21X1 OAI21X1_588 ( .A(_4552_), .B(decoded_imm_0_), .C(_4539__bF_buf1), .Y(_5851_) );
OAI22X1 OAI22X1_12 ( .A(_5142_), .B(_4539__bF_buf0), .C(_5850_), .D(_5851_), .Y(_82__0_) );
NOR2X1 NOR2X1_264 ( .A(_5849__bF_buf3), .B(_5488_), .Y(_5852_) );
OAI21X1 OAI21X1_589 ( .A(_4552_), .B(decoded_imm_1_), .C(_4539__bF_buf3), .Y(_5853_) );
OAI22X1 OAI22X1_13 ( .A(_5140__bF_buf3), .B(_4539__bF_buf2), .C(_5852_), .D(_5853_), .Y(_82__1_) );
NOR2X1 NOR2X1_265 ( .A(_5849__bF_buf2), .B(_5560_), .Y(_5854_) );
OAI21X1 OAI21X1_590 ( .A(_4552_), .B(decoded_imm_2_), .C(_4539__bF_buf1), .Y(_5855_) );
OAI22X1 OAI22X1_14 ( .A(_5131__bF_buf3), .B(_4539__bF_buf0), .C(_5854_), .D(_5855_), .Y(_82__2_) );
INVX1 INVX1_342 ( .A(_10728__3_bF_buf1_), .Y(_5856_) );
NOR2X1 NOR2X1_266 ( .A(_5849__bF_buf1), .B(_5629_), .Y(_5857_) );
OAI21X1 OAI21X1_591 ( .A(_4552_), .B(decoded_imm_3_), .C(_4539__bF_buf3), .Y(_5858_) );
OAI22X1 OAI22X1_15 ( .A(_5856__bF_buf4), .B(_4539__bF_buf2), .C(_5857_), .D(_5858_), .Y(_82__3_) );
INVX1 INVX1_343 ( .A(_10728__4_bF_buf1_), .Y(_5859_) );
NOR2X1 NOR2X1_267 ( .A(_5849__bF_buf0), .B(_5700_), .Y(_5860_) );
OAI21X1 OAI21X1_592 ( .A(_4552_), .B(decoded_imm_4_), .C(_4539__bF_buf1), .Y(_5861_) );
OAI22X1 OAI22X1_16 ( .A(_5859__bF_buf4), .B(_4539__bF_buf0), .C(_5860_), .D(_5861_), .Y(_82__4_) );
INVX1 INVX1_344 ( .A(_10728__5_), .Y(_5862_) );
NOR2X1 NOR2X1_268 ( .A(decoded_rs2_0_bF_buf22_), .B(cpuregs_0_[5]), .Y(_5863_) );
OAI21X1 OAI21X1_593 ( .A(_5362__bF_buf5), .B(cpuregs_1_[5]), .C(_5349__bF_buf7), .Y(_5864_) );
NOR2X1 NOR2X1_269 ( .A(cpuregs_3_[5]), .B(_5362__bF_buf4), .Y(_5865_) );
OAI21X1 OAI21X1_594 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_2_[5]), .C(decoded_rs2_1_bF_buf7_), .Y(_5866_) );
OAI22X1 OAI22X1_17 ( .A(_5865_), .B(_5866_), .C(_5864_), .D(_5863_), .Y(_5867_) );
NOR2X1 NOR2X1_270 ( .A(decoded_rs2_2_bF_buf0_), .B(_5867_), .Y(_5868_) );
NOR2X1 NOR2X1_271 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_4_[5]), .Y(_5869_) );
OAI21X1 OAI21X1_595 ( .A(_5362__bF_buf3), .B(cpuregs_5_[5]), .C(_5349__bF_buf6), .Y(_5870_) );
NOR2X1 NOR2X1_272 ( .A(cpuregs_7_[5]), .B(_5362__bF_buf2), .Y(_5871_) );
OAI21X1 OAI21X1_596 ( .A(cpuregs_6_[5]), .B(decoded_rs2_0_bF_buf19_), .C(decoded_rs2_1_bF_buf6_), .Y(_5872_) );
OAI22X1 OAI22X1_18 ( .A(_5871_), .B(_5872_), .C(_5870_), .D(_5869_), .Y(_5873_) );
OAI21X1 OAI21X1_597 ( .A(_5873_), .B(_5358__bF_buf11), .C(_5348__bF_buf1), .Y(_5874_) );
INVX1 INVX1_345 ( .A(cpuregs_9_[5]), .Y(_5875_) );
AOI21X1 AOI21X1_65 ( .A(decoded_rs2_0_bF_buf18_), .B(_5875_), .C(decoded_rs2_1_bF_buf5_), .Y(_5876_) );
OAI21X1 OAI21X1_598 ( .A(cpuregs_8_[5]), .B(decoded_rs2_0_bF_buf17_), .C(_5876_), .Y(_5877_) );
NOR2X1 NOR2X1_273 ( .A(cpuregs_11_[5]), .B(_5362__bF_buf1), .Y(_5878_) );
OAI21X1 OAI21X1_599 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_10_[5]), .C(decoded_rs2_1_bF_buf4_), .Y(_5879_) );
OAI21X1 OAI21X1_600 ( .A(_5878_), .B(_5879_), .C(_5877_), .Y(_5880_) );
NOR2X1 NOR2X1_274 ( .A(decoded_rs2_2_bF_buf8_), .B(_5880_), .Y(_5881_) );
NOR2X1 NOR2X1_275 ( .A(decoded_rs2_0_bF_buf15_), .B(cpuregs_12_[5]), .Y(_5882_) );
OAI21X1 OAI21X1_601 ( .A(_5362__bF_buf0), .B(cpuregs_13_[5]), .C(_5349__bF_buf5), .Y(_5883_) );
INVX1 INVX1_346 ( .A(cpuregs_14_[5]), .Y(_5884_) );
AOI21X1 AOI21X1_66 ( .A(_5362__bF_buf14), .B(_5884_), .C(_5349__bF_buf4), .Y(_5885_) );
OAI21X1 OAI21X1_602 ( .A(_5362__bF_buf13), .B(cpuregs_15_[5]), .C(_5885_), .Y(_5886_) );
OAI21X1 OAI21X1_603 ( .A(_5882_), .B(_5883_), .C(_5886_), .Y(_5887_) );
OAI21X1 OAI21X1_604 ( .A(_5887_), .B(_5358__bF_buf10), .C(decoded_rs2_3_bF_buf1_), .Y(_5888_) );
OAI22X1 OAI22X1_19 ( .A(_5868_), .B(_5874_), .C(_5888_), .D(_5881_), .Y(_5889_) );
OAI21X1 OAI21X1_605 ( .A(_5385_), .B(_5384_), .C(_4552_), .Y(_5890_) );
INVX1 INVX1_347 ( .A(cpuregs_26_[5]), .Y(_5891_) );
OAI21X1 OAI21X1_606 ( .A(_5891_), .B(decoded_rs2_0_bF_buf14_), .C(decoded_rs2_1_bF_buf3_), .Y(_5892_) );
AOI21X1 AOI21X1_67 ( .A(decoded_rs2_0_bF_buf13_), .B(cpuregs_27_[5]), .C(_5892_), .Y(_5893_) );
AND2X2 AND2X2_23 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_25_[5]), .Y(_5894_) );
INVX1 INVX1_348 ( .A(cpuregs_24_[5]), .Y(_5895_) );
OAI21X1 OAI21X1_607 ( .A(_5895_), .B(decoded_rs2_0_bF_buf11_), .C(_5349__bF_buf3), .Y(_5896_) );
OAI21X1 OAI21X1_608 ( .A(_5896_), .B(_5894_), .C(_5358__bF_buf9), .Y(_5897_) );
INVX1 INVX1_349 ( .A(cpuregs_28_[5]), .Y(_5898_) );
NAND2X1 NAND2X1_327 ( .A(decoded_rs2_0_bF_buf10_), .B(cpuregs_29_[5]), .Y(_5899_) );
OAI21X1 OAI21X1_609 ( .A(_5898_), .B(decoded_rs2_0_bF_buf9_), .C(_5899_), .Y(_5900_) );
INVX1 INVX1_350 ( .A(cpuregs_30_[5]), .Y(_5901_) );
NAND2X1 NAND2X1_328 ( .A(decoded_rs2_0_bF_buf8_), .B(cpuregs_31_[5]), .Y(_5902_) );
OAI21X1 OAI21X1_610 ( .A(_5901_), .B(decoded_rs2_0_bF_buf7_), .C(_5902_), .Y(_5903_) );
MUX2X1 MUX2X1_60 ( .A(_5903_), .B(_5900_), .S(decoded_rs2_1_bF_buf2_), .Y(_5904_) );
OAI22X1 OAI22X1_20 ( .A(_5897_), .B(_5893_), .C(_5904_), .D(_5358__bF_buf8), .Y(_5905_) );
INVX1 INVX1_351 ( .A(cpuregs_16_[5]), .Y(_5906_) );
NAND2X1 NAND2X1_329 ( .A(decoded_rs2_0_bF_buf6_), .B(cpuregs_17_[5]), .Y(_5907_) );
OAI21X1 OAI21X1_611 ( .A(_5906_), .B(decoded_rs2_0_bF_buf5_), .C(_5907_), .Y(_5908_) );
INVX1 INVX1_352 ( .A(cpuregs_18_[5]), .Y(_5909_) );
NAND2X1 NAND2X1_330 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_19_[5]), .Y(_5910_) );
OAI21X1 OAI21X1_612 ( .A(_5909_), .B(decoded_rs2_0_bF_buf3_), .C(_5910_), .Y(_5911_) );
MUX2X1 MUX2X1_61 ( .A(_5911_), .B(_5908_), .S(decoded_rs2_1_bF_buf1_), .Y(_5912_) );
NAND2X1 NAND2X1_331 ( .A(_5358__bF_buf7), .B(_5912_), .Y(_5913_) );
INVX1 INVX1_353 ( .A(cpuregs_20_[5]), .Y(_5914_) );
NAND2X1 NAND2X1_332 ( .A(decoded_rs2_0_bF_buf2_), .B(cpuregs_21_[5]), .Y(_5915_) );
OAI21X1 OAI21X1_613 ( .A(_5914_), .B(decoded_rs2_0_bF_buf1_), .C(_5915_), .Y(_5916_) );
INVX1 INVX1_354 ( .A(cpuregs_23_[5]), .Y(_5917_) );
NAND2X1 NAND2X1_333 ( .A(cpuregs_22_[5]), .B(_5362__bF_buf12), .Y(_5918_) );
OAI21X1 OAI21X1_614 ( .A(_5362__bF_buf11), .B(_5917_), .C(_5918_), .Y(_5919_) );
MUX2X1 MUX2X1_62 ( .A(_5919_), .B(_5916_), .S(decoded_rs2_1_bF_buf0_), .Y(_5920_) );
AOI21X1 AOI21X1_68 ( .A(decoded_rs2_2_bF_buf7_), .B(_5920_), .C(decoded_rs2_3_bF_buf0_), .Y(_5921_) );
AOI22X1 AOI22X1_12 ( .A(decoded_rs2_3_bF_buf6_), .B(_5905_), .C(_5921_), .D(_5913_), .Y(_5922_) );
AOI21X1 AOI21X1_69 ( .A(decoded_rs2_4_bF_buf0_), .B(_5922_), .C(_5890__bF_buf3), .Y(_5923_) );
OAI21X1 OAI21X1_615 ( .A(decoded_rs2_4_bF_buf7_), .B(_5889_), .C(_5923_), .Y(_5924_) );
AOI21X1 AOI21X1_70 ( .A(decoded_imm_5_), .B(_5849__bF_buf4), .C(_4540__bF_buf5), .Y(_5925_) );
AOI22X1 AOI22X1_13 ( .A(_5862_), .B(_4540__bF_buf4), .C(_5924_), .D(_5925_), .Y(_82__5_) );
INVX1 INVX1_355 ( .A(_10728__6_), .Y(_5926_) );
NOR2X1 NOR2X1_276 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_0_[6]), .Y(_5927_) );
OAI21X1 OAI21X1_616 ( .A(_5362__bF_buf10), .B(cpuregs_1_[6]), .C(_5349__bF_buf2), .Y(_5928_) );
NOR2X1 NOR2X1_277 ( .A(cpuregs_3_[6]), .B(_5362__bF_buf9), .Y(_5929_) );
OAI21X1 OAI21X1_617 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_2_[6]), .C(decoded_rs2_1_bF_buf45_), .Y(_5930_) );
OAI22X1 OAI22X1_21 ( .A(_5929_), .B(_5930_), .C(_5928_), .D(_5927_), .Y(_5931_) );
NOR2X1 NOR2X1_278 ( .A(decoded_rs2_2_bF_buf6_), .B(_5931_), .Y(_5932_) );
NOR2X1 NOR2X1_279 ( .A(decoded_rs2_0_bF_buf77_), .B(cpuregs_4_[6]), .Y(_5933_) );
OAI21X1 OAI21X1_618 ( .A(_5362__bF_buf8), .B(cpuregs_5_[6]), .C(_5349__bF_buf1), .Y(_5934_) );
NOR2X1 NOR2X1_280 ( .A(cpuregs_7_[6]), .B(_5362__bF_buf7), .Y(_5935_) );
OAI21X1 OAI21X1_619 ( .A(cpuregs_6_[6]), .B(decoded_rs2_0_bF_buf76_), .C(decoded_rs2_1_bF_buf44_), .Y(_5936_) );
OAI22X1 OAI22X1_22 ( .A(_5935_), .B(_5936_), .C(_5934_), .D(_5933_), .Y(_5937_) );
OAI21X1 OAI21X1_620 ( .A(_5937_), .B(_5358__bF_buf6), .C(_5348__bF_buf0), .Y(_5938_) );
INVX1 INVX1_356 ( .A(cpuregs_9_[6]), .Y(_5939_) );
AOI21X1 AOI21X1_71 ( .A(decoded_rs2_0_bF_buf75_), .B(_5939_), .C(decoded_rs2_1_bF_buf43_), .Y(_5940_) );
OAI21X1 OAI21X1_621 ( .A(cpuregs_8_[6]), .B(decoded_rs2_0_bF_buf74_), .C(_5940_), .Y(_5941_) );
INVX1 INVX1_357 ( .A(cpuregs_10_[6]), .Y(_5942_) );
AOI21X1 AOI21X1_72 ( .A(_5362__bF_buf6), .B(_5942_), .C(_5349__bF_buf0), .Y(_5943_) );
OAI21X1 OAI21X1_622 ( .A(_5362__bF_buf5), .B(cpuregs_11_[6]), .C(_5943_), .Y(_5944_) );
AOI21X1 AOI21X1_73 ( .A(_5941_), .B(_5944_), .C(decoded_rs2_2_bF_buf5_), .Y(_5945_) );
NOR2X1 NOR2X1_281 ( .A(decoded_rs2_0_bF_buf73_), .B(cpuregs_12_[6]), .Y(_5946_) );
OAI21X1 OAI21X1_623 ( .A(_5362__bF_buf4), .B(cpuregs_13_[6]), .C(_5349__bF_buf11), .Y(_5947_) );
INVX1 INVX1_358 ( .A(cpuregs_14_[6]), .Y(_5948_) );
AOI21X1 AOI21X1_74 ( .A(_5362__bF_buf3), .B(_5948_), .C(_5349__bF_buf10), .Y(_5949_) );
OAI21X1 OAI21X1_624 ( .A(_5362__bF_buf2), .B(cpuregs_15_[6]), .C(_5949_), .Y(_5950_) );
OAI21X1 OAI21X1_625 ( .A(_5946_), .B(_5947_), .C(_5950_), .Y(_5951_) );
AND2X2 AND2X2_24 ( .A(_5951_), .B(decoded_rs2_2_bF_buf4_), .Y(_5952_) );
OAI21X1 OAI21X1_626 ( .A(_5952_), .B(_5945_), .C(decoded_rs2_3_bF_buf5_), .Y(_5953_) );
OAI21X1 OAI21X1_627 ( .A(_5932_), .B(_5938_), .C(_5953_), .Y(_5954_) );
INVX1 INVX1_359 ( .A(cpuregs_26_[6]), .Y(_5955_) );
OAI21X1 OAI21X1_628 ( .A(_5955_), .B(decoded_rs2_0_bF_buf72_), .C(decoded_rs2_1_bF_buf42_), .Y(_5956_) );
AOI21X1 AOI21X1_75 ( .A(decoded_rs2_0_bF_buf71_), .B(cpuregs_27_[6]), .C(_5956_), .Y(_5957_) );
AND2X2 AND2X2_25 ( .A(decoded_rs2_0_bF_buf70_), .B(cpuregs_25_[6]), .Y(_5958_) );
INVX1 INVX1_360 ( .A(cpuregs_24_[6]), .Y(_5959_) );
OAI21X1 OAI21X1_629 ( .A(_5959_), .B(decoded_rs2_0_bF_buf69_), .C(_5349__bF_buf9), .Y(_5960_) );
OAI21X1 OAI21X1_630 ( .A(_5960_), .B(_5958_), .C(_5358__bF_buf5), .Y(_5961_) );
INVX1 INVX1_361 ( .A(cpuregs_28_[6]), .Y(_5962_) );
NAND2X1 NAND2X1_334 ( .A(decoded_rs2_0_bF_buf68_), .B(cpuregs_29_[6]), .Y(_5963_) );
OAI21X1 OAI21X1_631 ( .A(_5962_), .B(decoded_rs2_0_bF_buf67_), .C(_5963_), .Y(_5964_) );
INVX1 INVX1_362 ( .A(cpuregs_30_[6]), .Y(_5965_) );
NAND2X1 NAND2X1_335 ( .A(decoded_rs2_0_bF_buf66_), .B(cpuregs_31_[6]), .Y(_5966_) );
OAI21X1 OAI21X1_632 ( .A(_5965_), .B(decoded_rs2_0_bF_buf65_), .C(_5966_), .Y(_5967_) );
MUX2X1 MUX2X1_63 ( .A(_5967_), .B(_5964_), .S(decoded_rs2_1_bF_buf41_), .Y(_5968_) );
OAI22X1 OAI22X1_23 ( .A(_5961_), .B(_5957_), .C(_5968_), .D(_5358__bF_buf4), .Y(_5969_) );
INVX1 INVX1_363 ( .A(cpuregs_16_[6]), .Y(_5970_) );
NAND2X1 NAND2X1_336 ( .A(decoded_rs2_0_bF_buf64_), .B(cpuregs_17_[6]), .Y(_5971_) );
OAI21X1 OAI21X1_633 ( .A(_5970_), .B(decoded_rs2_0_bF_buf63_), .C(_5971_), .Y(_5972_) );
INVX1 INVX1_364 ( .A(cpuregs_18_[6]), .Y(_5973_) );
NAND2X1 NAND2X1_337 ( .A(decoded_rs2_0_bF_buf62_), .B(cpuregs_19_[6]), .Y(_5974_) );
OAI21X1 OAI21X1_634 ( .A(_5973_), .B(decoded_rs2_0_bF_buf61_), .C(_5974_), .Y(_5975_) );
MUX2X1 MUX2X1_64 ( .A(_5975_), .B(_5972_), .S(decoded_rs2_1_bF_buf40_), .Y(_5976_) );
NAND2X1 NAND2X1_338 ( .A(_5358__bF_buf3), .B(_5976_), .Y(_5977_) );
INVX1 INVX1_365 ( .A(cpuregs_20_[6]), .Y(_5978_) );
NAND2X1 NAND2X1_339 ( .A(decoded_rs2_0_bF_buf60_), .B(cpuregs_21_[6]), .Y(_5979_) );
OAI21X1 OAI21X1_635 ( .A(_5978_), .B(decoded_rs2_0_bF_buf59_), .C(_5979_), .Y(_5980_) );
INVX1 INVX1_366 ( .A(cpuregs_23_[6]), .Y(_5981_) );
NAND2X1 NAND2X1_340 ( .A(cpuregs_22_[6]), .B(_5362__bF_buf1), .Y(_5982_) );
OAI21X1 OAI21X1_636 ( .A(_5362__bF_buf0), .B(_5981_), .C(_5982_), .Y(_5983_) );
MUX2X1 MUX2X1_65 ( .A(_5983_), .B(_5980_), .S(decoded_rs2_1_bF_buf39_), .Y(_5984_) );
AOI21X1 AOI21X1_76 ( .A(decoded_rs2_2_bF_buf3_), .B(_5984_), .C(decoded_rs2_3_bF_buf4_), .Y(_5985_) );
AOI22X1 AOI22X1_14 ( .A(decoded_rs2_3_bF_buf3_), .B(_5969_), .C(_5985_), .D(_5977_), .Y(_5986_) );
AOI21X1 AOI21X1_77 ( .A(decoded_rs2_4_bF_buf6_), .B(_5986_), .C(_5890__bF_buf2), .Y(_5987_) );
OAI21X1 OAI21X1_637 ( .A(_5954_), .B(decoded_rs2_4_bF_buf5_), .C(_5987_), .Y(_5988_) );
AOI21X1 AOI21X1_78 ( .A(decoded_imm_6_), .B(_5849__bF_buf3), .C(_4540__bF_buf3), .Y(_5989_) );
AOI22X1 AOI22X1_15 ( .A(_5926_), .B(_4540__bF_buf2), .C(_5988_), .D(_5989_), .Y(_82__6_) );
INVX1 INVX1_367 ( .A(_10728__7_), .Y(_5990_) );
INVX1 INVX1_368 ( .A(cpuregs_9_[7]), .Y(_5991_) );
AOI21X1 AOI21X1_79 ( .A(decoded_rs2_0_bF_buf58_), .B(_5991_), .C(decoded_rs2_1_bF_buf38_), .Y(_5992_) );
OAI21X1 OAI21X1_638 ( .A(cpuregs_8_[7]), .B(decoded_rs2_0_bF_buf57_), .C(_5992_), .Y(_5993_) );
NOR2X1 NOR2X1_282 ( .A(cpuregs_11_[7]), .B(_5362__bF_buf14), .Y(_5994_) );
OAI21X1 OAI21X1_639 ( .A(decoded_rs2_0_bF_buf56_), .B(cpuregs_10_[7]), .C(decoded_rs2_1_bF_buf37_), .Y(_5995_) );
OAI21X1 OAI21X1_640 ( .A(_5994_), .B(_5995_), .C(_5993_), .Y(_5996_) );
NOR2X1 NOR2X1_283 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_12_[7]), .Y(_5997_) );
OAI21X1 OAI21X1_641 ( .A(_5362__bF_buf13), .B(cpuregs_13_[7]), .C(_5349__bF_buf8), .Y(_5998_) );
NOR2X1 NOR2X1_284 ( .A(cpuregs_15_[7]), .B(_5362__bF_buf12), .Y(_5999_) );
OAI21X1 OAI21X1_642 ( .A(decoded_rs2_0_bF_buf54_), .B(cpuregs_14_[7]), .C(decoded_rs2_1_bF_buf36_), .Y(_6000_) );
OAI22X1 OAI22X1_24 ( .A(_5999_), .B(_6000_), .C(_5998_), .D(_5997_), .Y(_6001_) );
MUX2X1 MUX2X1_66 ( .A(_5996_), .B(_6001_), .S(_5358__bF_buf2), .Y(_6002_) );
NOR2X1 NOR2X1_285 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_4_[7]), .Y(_6003_) );
OAI21X1 OAI21X1_643 ( .A(_5362__bF_buf11), .B(cpuregs_5_[7]), .C(_5349__bF_buf7), .Y(_6004_) );
NOR2X1 NOR2X1_286 ( .A(cpuregs_7_[7]), .B(_5362__bF_buf10), .Y(_6005_) );
OAI21X1 OAI21X1_644 ( .A(cpuregs_6_[7]), .B(decoded_rs2_0_bF_buf52_), .C(decoded_rs2_1_bF_buf35_), .Y(_6006_) );
OAI22X1 OAI22X1_25 ( .A(_6005_), .B(_6006_), .C(_6004_), .D(_6003_), .Y(_6007_) );
NOR2X1 NOR2X1_287 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_0_[7]), .Y(_6008_) );
OAI21X1 OAI21X1_645 ( .A(_5362__bF_buf9), .B(cpuregs_1_[7]), .C(_5349__bF_buf6), .Y(_6009_) );
NOR2X1 NOR2X1_288 ( .A(cpuregs_3_[7]), .B(_5362__bF_buf8), .Y(_6010_) );
OAI21X1 OAI21X1_646 ( .A(decoded_rs2_0_bF_buf50_), .B(cpuregs_2_[7]), .C(decoded_rs2_1_bF_buf34_), .Y(_6011_) );
OAI22X1 OAI22X1_26 ( .A(_6010_), .B(_6011_), .C(_6009_), .D(_6008_), .Y(_6012_) );
MUX2X1 MUX2X1_67 ( .A(_6012_), .B(_6007_), .S(_5358__bF_buf1), .Y(_6013_) );
MUX2X1 MUX2X1_68 ( .A(_6002_), .B(_6013_), .S(decoded_rs2_3_bF_buf2_), .Y(_6014_) );
INVX1 INVX1_369 ( .A(cpuregs_16_[7]), .Y(_6015_) );
NAND2X1 NAND2X1_341 ( .A(decoded_rs2_0_bF_buf49_), .B(cpuregs_17_[7]), .Y(_6016_) );
OAI21X1 OAI21X1_647 ( .A(_6015_), .B(decoded_rs2_0_bF_buf48_), .C(_6016_), .Y(_6017_) );
INVX1 INVX1_370 ( .A(cpuregs_18_[7]), .Y(_6018_) );
NAND2X1 NAND2X1_342 ( .A(decoded_rs2_0_bF_buf47_), .B(cpuregs_19_[7]), .Y(_6019_) );
OAI21X1 OAI21X1_648 ( .A(_6018_), .B(decoded_rs2_0_bF_buf46_), .C(_6019_), .Y(_6020_) );
MUX2X1 MUX2X1_69 ( .A(_6020_), .B(_6017_), .S(decoded_rs2_1_bF_buf33_), .Y(_6021_) );
NOR2X1 NOR2X1_289 ( .A(decoded_rs2_2_bF_buf2_), .B(_6021_), .Y(_6022_) );
INVX1 INVX1_371 ( .A(cpuregs_20_[7]), .Y(_6023_) );
NAND2X1 NAND2X1_343 ( .A(decoded_rs2_0_bF_buf45_), .B(cpuregs_21_[7]), .Y(_6024_) );
OAI21X1 OAI21X1_649 ( .A(_6023_), .B(decoded_rs2_0_bF_buf44_), .C(_6024_), .Y(_6025_) );
INVX1 INVX1_372 ( .A(cpuregs_23_[7]), .Y(_6026_) );
NAND2X1 NAND2X1_344 ( .A(cpuregs_22_[7]), .B(_5362__bF_buf7), .Y(_6027_) );
OAI21X1 OAI21X1_650 ( .A(_5362__bF_buf6), .B(_6026_), .C(_6027_), .Y(_6028_) );
MUX2X1 MUX2X1_70 ( .A(_6028_), .B(_6025_), .S(decoded_rs2_1_bF_buf32_), .Y(_6029_) );
NOR2X1 NOR2X1_290 ( .A(_5358__bF_buf0), .B(_6029_), .Y(_6030_) );
OAI21X1 OAI21X1_651 ( .A(_6030_), .B(_6022_), .C(_5348__bF_buf5), .Y(_6031_) );
INVX1 INVX1_373 ( .A(cpuregs_25_[7]), .Y(_6032_) );
AOI21X1 AOI21X1_80 ( .A(decoded_rs2_0_bF_buf43_), .B(_6032_), .C(decoded_rs2_1_bF_buf31_), .Y(_6033_) );
OAI21X1 OAI21X1_652 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_24_[7]), .C(_6033_), .Y(_6034_) );
NOR2X1 NOR2X1_291 ( .A(cpuregs_27_[7]), .B(_5362__bF_buf5), .Y(_6035_) );
OAI21X1 OAI21X1_653 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_26_[7]), .C(decoded_rs2_1_bF_buf30_), .Y(_6036_) );
OAI21X1 OAI21X1_654 ( .A(_6035_), .B(_6036_), .C(_6034_), .Y(_6037_) );
NOR2X1 NOR2X1_292 ( .A(decoded_rs2_2_bF_buf1_), .B(_6037_), .Y(_6038_) );
NOR2X1 NOR2X1_293 ( .A(decoded_rs2_0_bF_buf40_), .B(cpuregs_28_[7]), .Y(_6039_) );
OAI21X1 OAI21X1_655 ( .A(_5362__bF_buf4), .B(cpuregs_29_[7]), .C(_5349__bF_buf5), .Y(_6040_) );
INVX1 INVX1_374 ( .A(cpuregs_30_[7]), .Y(_6041_) );
AOI21X1 AOI21X1_81 ( .A(_5362__bF_buf3), .B(_6041_), .C(_5349__bF_buf4), .Y(_6042_) );
OAI21X1 OAI21X1_656 ( .A(_5362__bF_buf2), .B(cpuregs_31_[7]), .C(_6042_), .Y(_6043_) );
OAI21X1 OAI21X1_657 ( .A(_6039_), .B(_6040_), .C(_6043_), .Y(_6044_) );
OAI21X1 OAI21X1_658 ( .A(_6044_), .B(_5358__bF_buf12), .C(decoded_rs2_3_bF_buf1_), .Y(_6045_) );
OAI21X1 OAI21X1_659 ( .A(_6038_), .B(_6045_), .C(_6031_), .Y(_6046_) );
NOR2X1 NOR2X1_294 ( .A(_5347_), .B(_6046_), .Y(_6047_) );
NOR2X1 NOR2X1_295 ( .A(_5890__bF_buf1), .B(_6047_), .Y(_6048_) );
OAI21X1 OAI21X1_660 ( .A(decoded_rs2_4_bF_buf4_), .B(_6014_), .C(_6048_), .Y(_6049_) );
AOI21X1 AOI21X1_82 ( .A(decoded_imm_7_), .B(_5849__bF_buf2), .C(_4540__bF_buf1), .Y(_6050_) );
AOI22X1 AOI22X1_16 ( .A(_5990_), .B(_4540__bF_buf0), .C(_6049_), .D(_6050_), .Y(_82__7_) );
INVX1 INVX1_375 ( .A(_10735__8_), .Y(_6051_) );
NOR2X1 NOR2X1_296 ( .A(decoded_rs2_0_bF_buf39_), .B(cpuregs_0_[8]), .Y(_6052_) );
OAI21X1 OAI21X1_661 ( .A(_5362__bF_buf1), .B(cpuregs_1_[8]), .C(_5349__bF_buf3), .Y(_6053_) );
NOR2X1 NOR2X1_297 ( .A(cpuregs_3_[8]), .B(_5362__bF_buf0), .Y(_6054_) );
OAI21X1 OAI21X1_662 ( .A(decoded_rs2_0_bF_buf38_), .B(cpuregs_2_[8]), .C(decoded_rs2_1_bF_buf29_), .Y(_6055_) );
OAI22X1 OAI22X1_27 ( .A(_6054_), .B(_6055_), .C(_6053_), .D(_6052_), .Y(_6056_) );
NOR2X1 NOR2X1_298 ( .A(decoded_rs2_2_bF_buf0_), .B(_6056_), .Y(_6057_) );
NOR2X1 NOR2X1_299 ( .A(decoded_rs2_0_bF_buf37_), .B(cpuregs_4_[8]), .Y(_6058_) );
OAI21X1 OAI21X1_663 ( .A(_5362__bF_buf14), .B(cpuregs_5_[8]), .C(_5349__bF_buf2), .Y(_6059_) );
NOR2X1 NOR2X1_300 ( .A(cpuregs_7_[8]), .B(_5362__bF_buf13), .Y(_6060_) );
OAI21X1 OAI21X1_664 ( .A(cpuregs_6_[8]), .B(decoded_rs2_0_bF_buf36_), .C(decoded_rs2_1_bF_buf28_), .Y(_6061_) );
OAI22X1 OAI22X1_28 ( .A(_6060_), .B(_6061_), .C(_6059_), .D(_6058_), .Y(_6062_) );
OAI21X1 OAI21X1_665 ( .A(_6062_), .B(_5358__bF_buf11), .C(_5348__bF_buf4), .Y(_6063_) );
NOR2X1 NOR2X1_301 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_12_[8]), .Y(_6064_) );
OAI21X1 OAI21X1_666 ( .A(_5362__bF_buf12), .B(cpuregs_13_[8]), .C(_5349__bF_buf1), .Y(_6065_) );
NOR2X1 NOR2X1_302 ( .A(cpuregs_15_[8]), .B(_5362__bF_buf11), .Y(_6066_) );
OAI21X1 OAI21X1_667 ( .A(decoded_rs2_0_bF_buf34_), .B(cpuregs_14_[8]), .C(decoded_rs2_1_bF_buf27_), .Y(_6067_) );
OAI22X1 OAI22X1_29 ( .A(_6066_), .B(_6067_), .C(_6065_), .D(_6064_), .Y(_6068_) );
NOR2X1 NOR2X1_303 ( .A(_5358__bF_buf10), .B(_6068_), .Y(_6069_) );
INVX1 INVX1_376 ( .A(cpuregs_9_[8]), .Y(_6070_) );
AOI21X1 AOI21X1_83 ( .A(decoded_rs2_0_bF_buf33_), .B(_6070_), .C(decoded_rs2_1_bF_buf26_), .Y(_6071_) );
OAI21X1 OAI21X1_668 ( .A(cpuregs_8_[8]), .B(decoded_rs2_0_bF_buf32_), .C(_6071_), .Y(_6072_) );
NOR2X1 NOR2X1_304 ( .A(cpuregs_11_[8]), .B(_5362__bF_buf10), .Y(_6073_) );
OAI21X1 OAI21X1_669 ( .A(decoded_rs2_0_bF_buf31_), .B(cpuregs_10_[8]), .C(decoded_rs2_1_bF_buf25_), .Y(_6074_) );
OAI21X1 OAI21X1_670 ( .A(_6073_), .B(_6074_), .C(_6072_), .Y(_6075_) );
OAI21X1 OAI21X1_671 ( .A(_6075_), .B(decoded_rs2_2_bF_buf8_), .C(decoded_rs2_3_bF_buf0_), .Y(_6076_) );
OAI22X1 OAI22X1_30 ( .A(_6057_), .B(_6063_), .C(_6076_), .D(_6069_), .Y(_6077_) );
INVX1 INVX1_377 ( .A(cpuregs_26_[8]), .Y(_6078_) );
OAI21X1 OAI21X1_672 ( .A(_6078_), .B(decoded_rs2_0_bF_buf30_), .C(decoded_rs2_1_bF_buf24_), .Y(_6079_) );
AOI21X1 AOI21X1_84 ( .A(decoded_rs2_0_bF_buf29_), .B(cpuregs_27_[8]), .C(_6079_), .Y(_6080_) );
AND2X2 AND2X2_26 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_25_[8]), .Y(_6081_) );
INVX1 INVX1_378 ( .A(cpuregs_24_[8]), .Y(_6082_) );
OAI21X1 OAI21X1_673 ( .A(_6082_), .B(decoded_rs2_0_bF_buf27_), .C(_5349__bF_buf0), .Y(_6083_) );
OAI21X1 OAI21X1_674 ( .A(_6083_), .B(_6081_), .C(_5358__bF_buf9), .Y(_6084_) );
INVX1 INVX1_379 ( .A(cpuregs_28_[8]), .Y(_6085_) );
NAND2X1 NAND2X1_345 ( .A(decoded_rs2_0_bF_buf26_), .B(cpuregs_29_[8]), .Y(_6086_) );
OAI21X1 OAI21X1_675 ( .A(_6085_), .B(decoded_rs2_0_bF_buf25_), .C(_6086_), .Y(_6087_) );
INVX1 INVX1_380 ( .A(cpuregs_30_[8]), .Y(_6088_) );
NAND2X1 NAND2X1_346 ( .A(decoded_rs2_0_bF_buf24_), .B(cpuregs_31_[8]), .Y(_6089_) );
OAI21X1 OAI21X1_676 ( .A(_6088_), .B(decoded_rs2_0_bF_buf23_), .C(_6089_), .Y(_6090_) );
MUX2X1 MUX2X1_71 ( .A(_6090_), .B(_6087_), .S(decoded_rs2_1_bF_buf23_), .Y(_6091_) );
OAI22X1 OAI22X1_31 ( .A(_6084_), .B(_6080_), .C(_6091_), .D(_5358__bF_buf8), .Y(_6092_) );
INVX1 INVX1_381 ( .A(cpuregs_16_[8]), .Y(_6093_) );
NAND2X1 NAND2X1_347 ( .A(decoded_rs2_0_bF_buf22_), .B(cpuregs_17_[8]), .Y(_6094_) );
OAI21X1 OAI21X1_677 ( .A(_6093_), .B(decoded_rs2_0_bF_buf21_), .C(_6094_), .Y(_6095_) );
INVX1 INVX1_382 ( .A(cpuregs_18_[8]), .Y(_6096_) );
NAND2X1 NAND2X1_348 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_19_[8]), .Y(_6097_) );
OAI21X1 OAI21X1_678 ( .A(_6096_), .B(decoded_rs2_0_bF_buf19_), .C(_6097_), .Y(_6098_) );
MUX2X1 MUX2X1_72 ( .A(_6098_), .B(_6095_), .S(decoded_rs2_1_bF_buf22_), .Y(_6099_) );
NAND2X1 NAND2X1_349 ( .A(_5358__bF_buf7), .B(_6099_), .Y(_6100_) );
INVX1 INVX1_383 ( .A(cpuregs_20_[8]), .Y(_6101_) );
NAND2X1 NAND2X1_350 ( .A(decoded_rs2_0_bF_buf18_), .B(cpuregs_21_[8]), .Y(_6102_) );
OAI21X1 OAI21X1_679 ( .A(_6101_), .B(decoded_rs2_0_bF_buf17_), .C(_6102_), .Y(_6103_) );
INVX1 INVX1_384 ( .A(cpuregs_23_[8]), .Y(_6104_) );
NAND2X1 NAND2X1_351 ( .A(cpuregs_22_[8]), .B(_5362__bF_buf9), .Y(_6105_) );
OAI21X1 OAI21X1_680 ( .A(_5362__bF_buf8), .B(_6104_), .C(_6105_), .Y(_6106_) );
MUX2X1 MUX2X1_73 ( .A(_6106_), .B(_6103_), .S(decoded_rs2_1_bF_buf21_), .Y(_6107_) );
AOI21X1 AOI21X1_85 ( .A(decoded_rs2_2_bF_buf7_), .B(_6107_), .C(decoded_rs2_3_bF_buf6_), .Y(_6108_) );
AOI22X1 AOI22X1_17 ( .A(decoded_rs2_3_bF_buf5_), .B(_6092_), .C(_6108_), .D(_6100_), .Y(_6109_) );
AOI21X1 AOI21X1_86 ( .A(decoded_rs2_4_bF_buf3_), .B(_6109_), .C(_5890__bF_buf0), .Y(_6110_) );
OAI21X1 OAI21X1_681 ( .A(decoded_rs2_4_bF_buf2_), .B(_6077_), .C(_6110_), .Y(_6111_) );
AOI21X1 AOI21X1_87 ( .A(decoded_imm_8_), .B(_5849__bF_buf1), .C(_4540__bF_buf6), .Y(_6112_) );
AOI22X1 AOI22X1_18 ( .A(_6051_), .B(_4540__bF_buf5), .C(_6111_), .D(_6112_), .Y(_82__8_) );
INVX1 INVX1_385 ( .A(cpuregs_0_[9]), .Y(_6113_) );
NAND2X1 NAND2X1_352 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_1_[9]), .Y(_6114_) );
OAI21X1 OAI21X1_682 ( .A(_6113_), .B(decoded_rs2_0_bF_buf15_), .C(_6114_), .Y(_6115_) );
INVX1 INVX1_386 ( .A(cpuregs_2_[9]), .Y(_6116_) );
NAND2X1 NAND2X1_353 ( .A(decoded_rs2_0_bF_buf14_), .B(cpuregs_3_[9]), .Y(_6117_) );
OAI21X1 OAI21X1_683 ( .A(_6116_), .B(decoded_rs2_0_bF_buf13_), .C(_6117_), .Y(_6118_) );
MUX2X1 MUX2X1_74 ( .A(_6118_), .B(_6115_), .S(decoded_rs2_1_bF_buf20_), .Y(_6119_) );
NAND2X1 NAND2X1_354 ( .A(_5358__bF_buf6), .B(_6119_), .Y(_6120_) );
NOR2X1 NOR2X1_305 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_4_[9]), .Y(_6121_) );
OAI21X1 OAI21X1_684 ( .A(_5362__bF_buf7), .B(cpuregs_5_[9]), .C(_5349__bF_buf11), .Y(_6122_) );
NOR2X1 NOR2X1_306 ( .A(cpuregs_7_[9]), .B(_5362__bF_buf6), .Y(_6123_) );
OAI21X1 OAI21X1_685 ( .A(cpuregs_6_[9]), .B(decoded_rs2_0_bF_buf11_), .C(decoded_rs2_1_bF_buf19_), .Y(_6124_) );
OAI22X1 OAI22X1_32 ( .A(_6123_), .B(_6124_), .C(_6122_), .D(_6121_), .Y(_6125_) );
OAI21X1 OAI21X1_686 ( .A(_5358__bF_buf5), .B(_6125_), .C(_6120_), .Y(_6126_) );
INVX1 INVX1_387 ( .A(cpuregs_9_[9]), .Y(_6127_) );
AOI21X1 AOI21X1_88 ( .A(decoded_rs2_0_bF_buf10_), .B(_6127_), .C(decoded_rs2_1_bF_buf18_), .Y(_6128_) );
OAI21X1 OAI21X1_687 ( .A(cpuregs_8_[9]), .B(decoded_rs2_0_bF_buf9_), .C(_6128_), .Y(_6129_) );
NOR2X1 NOR2X1_307 ( .A(cpuregs_11_[9]), .B(_5362__bF_buf5), .Y(_6130_) );
OAI21X1 OAI21X1_688 ( .A(decoded_rs2_0_bF_buf8_), .B(cpuregs_10_[9]), .C(decoded_rs2_1_bF_buf17_), .Y(_6131_) );
OAI21X1 OAI21X1_689 ( .A(_6130_), .B(_6131_), .C(_6129_), .Y(_6132_) );
NOR2X1 NOR2X1_308 ( .A(decoded_rs2_2_bF_buf6_), .B(_6132_), .Y(_6133_) );
INVX1 INVX1_388 ( .A(cpuregs_13_[9]), .Y(_6134_) );
AOI21X1 AOI21X1_89 ( .A(decoded_rs2_0_bF_buf7_), .B(_6134_), .C(decoded_rs2_1_bF_buf16_), .Y(_6135_) );
OAI21X1 OAI21X1_690 ( .A(decoded_rs2_0_bF_buf6_), .B(cpuregs_12_[9]), .C(_6135_), .Y(_6136_) );
NOR2X1 NOR2X1_309 ( .A(cpuregs_15_[9]), .B(_5362__bF_buf4), .Y(_6137_) );
OAI21X1 OAI21X1_691 ( .A(decoded_rs2_0_bF_buf5_), .B(cpuregs_14_[9]), .C(decoded_rs2_1_bF_buf15_), .Y(_6138_) );
OAI21X1 OAI21X1_692 ( .A(_6137_), .B(_6138_), .C(_6136_), .Y(_6139_) );
OAI21X1 OAI21X1_693 ( .A(_6139_), .B(_5358__bF_buf4), .C(decoded_rs2_3_bF_buf4_), .Y(_6140_) );
OAI22X1 OAI22X1_33 ( .A(_6126_), .B(decoded_rs2_3_bF_buf3_), .C(_6133_), .D(_6140_), .Y(_6141_) );
INVX1 INVX1_389 ( .A(cpuregs_24_[9]), .Y(_6142_) );
NAND2X1 NAND2X1_355 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_25_[9]), .Y(_6143_) );
OAI21X1 OAI21X1_694 ( .A(_6142_), .B(decoded_rs2_0_bF_buf3_), .C(_6143_), .Y(_6144_) );
INVX1 INVX1_390 ( .A(cpuregs_27_[9]), .Y(_6145_) );
OAI21X1 OAI21X1_695 ( .A(decoded_rs2_0_bF_buf2_), .B(cpuregs_26_[9]), .C(decoded_rs2_1_bF_buf14_), .Y(_6146_) );
AOI21X1 AOI21X1_90 ( .A(decoded_rs2_0_bF_buf1_), .B(_6145_), .C(_6146_), .Y(_6147_) );
AOI21X1 AOI21X1_91 ( .A(_5349__bF_buf10), .B(_6144_), .C(_6147_), .Y(_6148_) );
INVX1 INVX1_391 ( .A(cpuregs_29_[9]), .Y(_6149_) );
NAND2X1 NAND2X1_356 ( .A(cpuregs_28_[9]), .B(_5362__bF_buf3), .Y(_6150_) );
OAI21X1 OAI21X1_696 ( .A(_5362__bF_buf2), .B(_6149_), .C(_6150_), .Y(_6151_) );
INVX1 INVX1_392 ( .A(cpuregs_31_[9]), .Y(_6152_) );
OAI21X1 OAI21X1_697 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_30_[9]), .C(decoded_rs2_1_bF_buf13_), .Y(_6153_) );
AOI21X1 AOI21X1_92 ( .A(decoded_rs2_0_bF_buf78_), .B(_6152_), .C(_6153_), .Y(_6154_) );
AOI21X1 AOI21X1_93 ( .A(_5349__bF_buf9), .B(_6151_), .C(_6154_), .Y(_6155_) );
MUX2X1 MUX2X1_75 ( .A(_6155_), .B(_6148_), .S(decoded_rs2_2_bF_buf5_), .Y(_6156_) );
INVX1 INVX1_393 ( .A(cpuregs_17_[9]), .Y(_6157_) );
NAND2X1 NAND2X1_357 ( .A(cpuregs_16_[9]), .B(_5362__bF_buf1), .Y(_6158_) );
OAI21X1 OAI21X1_698 ( .A(_5362__bF_buf0), .B(_6157_), .C(_6158_), .Y(_6159_) );
INVX1 INVX1_394 ( .A(cpuregs_19_[9]), .Y(_6160_) );
OAI21X1 OAI21X1_699 ( .A(decoded_rs2_0_bF_buf77_), .B(cpuregs_18_[9]), .C(decoded_rs2_1_bF_buf12_), .Y(_6161_) );
AOI21X1 AOI21X1_94 ( .A(decoded_rs2_0_bF_buf76_), .B(_6160_), .C(_6161_), .Y(_6162_) );
AOI21X1 AOI21X1_95 ( .A(_5349__bF_buf8), .B(_6159_), .C(_6162_), .Y(_6163_) );
NAND2X1 NAND2X1_358 ( .A(_5358__bF_buf3), .B(_6163_), .Y(_6164_) );
INVX1 INVX1_395 ( .A(cpuregs_20_[9]), .Y(_6165_) );
NAND2X1 NAND2X1_359 ( .A(decoded_rs2_0_bF_buf75_), .B(cpuregs_21_[9]), .Y(_6166_) );
OAI21X1 OAI21X1_700 ( .A(_6165_), .B(decoded_rs2_0_bF_buf74_), .C(_6166_), .Y(_6167_) );
INVX1 INVX1_396 ( .A(cpuregs_22_[9]), .Y(_6168_) );
NAND2X1 NAND2X1_360 ( .A(decoded_rs2_0_bF_buf73_), .B(cpuregs_23_[9]), .Y(_6169_) );
OAI21X1 OAI21X1_701 ( .A(_6168_), .B(decoded_rs2_0_bF_buf72_), .C(_6169_), .Y(_6170_) );
MUX2X1 MUX2X1_76 ( .A(_6170_), .B(_6167_), .S(decoded_rs2_1_bF_buf11_), .Y(_6171_) );
AOI21X1 AOI21X1_96 ( .A(decoded_rs2_2_bF_buf4_), .B(_6171_), .C(decoded_rs2_3_bF_buf2_), .Y(_6172_) );
AOI22X1 AOI22X1_19 ( .A(_6172_), .B(_6164_), .C(decoded_rs2_3_bF_buf1_), .D(_6156_), .Y(_6173_) );
AOI21X1 AOI21X1_97 ( .A(decoded_rs2_4_bF_buf1_), .B(_6173_), .C(_5890__bF_buf3), .Y(_6174_) );
OAI21X1 OAI21X1_702 ( .A(decoded_rs2_4_bF_buf0_), .B(_6141_), .C(_6174_), .Y(_6175_) );
AOI21X1 AOI21X1_98 ( .A(decoded_imm_9_), .B(_5849__bF_buf0), .C(_4540__bF_buf4), .Y(_6176_) );
AOI22X1 AOI22X1_20 ( .A(_5108_), .B(_4540__bF_buf3), .C(_6175_), .D(_6176_), .Y(_82__9_) );
INVX1 INVX1_397 ( .A(cpuregs_9_[10]), .Y(_6177_) );
AOI21X1 AOI21X1_99 ( .A(decoded_rs2_0_bF_buf71_), .B(_6177_), .C(decoded_rs2_1_bF_buf10_), .Y(_6178_) );
OAI21X1 OAI21X1_703 ( .A(cpuregs_8_[10]), .B(decoded_rs2_0_bF_buf70_), .C(_6178_), .Y(_6179_) );
NOR2X1 NOR2X1_310 ( .A(cpuregs_11_[10]), .B(_5362__bF_buf14), .Y(_6180_) );
OAI21X1 OAI21X1_704 ( .A(decoded_rs2_0_bF_buf69_), .B(cpuregs_10_[10]), .C(decoded_rs2_1_bF_buf9_), .Y(_6181_) );
OAI21X1 OAI21X1_705 ( .A(_6180_), .B(_6181_), .C(_6179_), .Y(_6182_) );
NOR2X1 NOR2X1_311 ( .A(decoded_rs2_0_bF_buf68_), .B(cpuregs_12_[10]), .Y(_6183_) );
OAI21X1 OAI21X1_706 ( .A(_5362__bF_buf13), .B(cpuregs_13_[10]), .C(_5349__bF_buf7), .Y(_6184_) );
NOR2X1 NOR2X1_312 ( .A(cpuregs_15_[10]), .B(_5362__bF_buf12), .Y(_6185_) );
OAI21X1 OAI21X1_707 ( .A(decoded_rs2_0_bF_buf67_), .B(cpuregs_14_[10]), .C(decoded_rs2_1_bF_buf8_), .Y(_6186_) );
OAI22X1 OAI22X1_34 ( .A(_6185_), .B(_6186_), .C(_6184_), .D(_6183_), .Y(_6187_) );
MUX2X1 MUX2X1_77 ( .A(_6182_), .B(_6187_), .S(_5358__bF_buf2), .Y(_6188_) );
NOR2X1 NOR2X1_313 ( .A(decoded_rs2_0_bF_buf66_), .B(cpuregs_4_[10]), .Y(_6189_) );
OAI21X1 OAI21X1_708 ( .A(_5362__bF_buf11), .B(cpuregs_5_[10]), .C(_5349__bF_buf6), .Y(_6190_) );
NOR2X1 NOR2X1_314 ( .A(cpuregs_7_[10]), .B(_5362__bF_buf10), .Y(_6191_) );
OAI21X1 OAI21X1_709 ( .A(cpuregs_6_[10]), .B(decoded_rs2_0_bF_buf65_), .C(decoded_rs2_1_bF_buf7_), .Y(_6192_) );
OAI22X1 OAI22X1_35 ( .A(_6191_), .B(_6192_), .C(_6190_), .D(_6189_), .Y(_6193_) );
NOR2X1 NOR2X1_315 ( .A(decoded_rs2_0_bF_buf64_), .B(cpuregs_0_[10]), .Y(_6194_) );
OAI21X1 OAI21X1_710 ( .A(_5362__bF_buf9), .B(cpuregs_1_[10]), .C(_5349__bF_buf5), .Y(_6195_) );
NOR2X1 NOR2X1_316 ( .A(cpuregs_3_[10]), .B(_5362__bF_buf8), .Y(_6196_) );
OAI21X1 OAI21X1_711 ( .A(decoded_rs2_0_bF_buf63_), .B(cpuregs_2_[10]), .C(decoded_rs2_1_bF_buf6_), .Y(_6197_) );
OAI22X1 OAI22X1_36 ( .A(_6196_), .B(_6197_), .C(_6195_), .D(_6194_), .Y(_6198_) );
MUX2X1 MUX2X1_78 ( .A(_6198_), .B(_6193_), .S(_5358__bF_buf1), .Y(_6199_) );
MUX2X1 MUX2X1_79 ( .A(_6188_), .B(_6199_), .S(decoded_rs2_3_bF_buf0_), .Y(_6200_) );
INVX1 INVX1_398 ( .A(cpuregs_17_[10]), .Y(_6201_) );
AOI21X1 AOI21X1_100 ( .A(decoded_rs2_0_bF_buf62_), .B(_6201_), .C(decoded_rs2_1_bF_buf5_), .Y(_6202_) );
OAI21X1 OAI21X1_712 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_16_[10]), .C(_6202_), .Y(_6203_) );
NOR2X1 NOR2X1_317 ( .A(cpuregs_19_[10]), .B(_5362__bF_buf7), .Y(_6204_) );
OAI21X1 OAI21X1_713 ( .A(decoded_rs2_0_bF_buf60_), .B(cpuregs_18_[10]), .C(decoded_rs2_1_bF_buf4_), .Y(_6205_) );
OAI21X1 OAI21X1_714 ( .A(_6204_), .B(_6205_), .C(_6203_), .Y(_6206_) );
INVX1 INVX1_399 ( .A(cpuregs_20_[10]), .Y(_6207_) );
NAND2X1 NAND2X1_361 ( .A(decoded_rs2_0_bF_buf59_), .B(cpuregs_21_[10]), .Y(_6208_) );
OAI21X1 OAI21X1_715 ( .A(_6207_), .B(decoded_rs2_0_bF_buf58_), .C(_6208_), .Y(_6209_) );
INVX1 INVX1_400 ( .A(cpuregs_23_[10]), .Y(_6210_) );
NAND2X1 NAND2X1_362 ( .A(cpuregs_22_[10]), .B(_5362__bF_buf6), .Y(_6211_) );
OAI21X1 OAI21X1_716 ( .A(_5362__bF_buf5), .B(_6210_), .C(_6211_), .Y(_6212_) );
MUX2X1 MUX2X1_80 ( .A(_6212_), .B(_6209_), .S(decoded_rs2_1_bF_buf3_), .Y(_6213_) );
NOR2X1 NOR2X1_318 ( .A(_5358__bF_buf0), .B(_6213_), .Y(_6214_) );
AOI21X1 AOI21X1_101 ( .A(_5358__bF_buf12), .B(_6206_), .C(_6214_), .Y(_6215_) );
NOR2X1 NOR2X1_319 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_24_[10]), .Y(_6216_) );
OAI21X1 OAI21X1_717 ( .A(_5362__bF_buf4), .B(cpuregs_25_[10]), .C(_5349__bF_buf4), .Y(_6217_) );
INVX1 INVX1_401 ( .A(cpuregs_26_[10]), .Y(_6218_) );
AOI21X1 AOI21X1_102 ( .A(_5362__bF_buf3), .B(_6218_), .C(_5349__bF_buf3), .Y(_6219_) );
OAI21X1 OAI21X1_718 ( .A(_5362__bF_buf2), .B(cpuregs_27_[10]), .C(_6219_), .Y(_6220_) );
OAI21X1 OAI21X1_719 ( .A(_6216_), .B(_6217_), .C(_6220_), .Y(_6221_) );
INVX1 INVX1_402 ( .A(cpuregs_28_[10]), .Y(_6222_) );
NAND2X1 NAND2X1_363 ( .A(decoded_rs2_0_bF_buf56_), .B(cpuregs_29_[10]), .Y(_6223_) );
OAI21X1 OAI21X1_720 ( .A(_6222_), .B(decoded_rs2_0_bF_buf55_), .C(_6223_), .Y(_6224_) );
INVX1 INVX1_403 ( .A(cpuregs_31_[10]), .Y(_6225_) );
OAI21X1 OAI21X1_721 ( .A(decoded_rs2_0_bF_buf54_), .B(cpuregs_30_[10]), .C(decoded_rs2_1_bF_buf2_), .Y(_6226_) );
AOI21X1 AOI21X1_103 ( .A(decoded_rs2_0_bF_buf53_), .B(_6225_), .C(_6226_), .Y(_6227_) );
AOI21X1 AOI21X1_104 ( .A(_5349__bF_buf2), .B(_6224_), .C(_6227_), .Y(_6228_) );
AOI21X1 AOI21X1_105 ( .A(decoded_rs2_2_bF_buf3_), .B(_6228_), .C(_5348__bF_buf3), .Y(_6229_) );
OAI21X1 OAI21X1_722 ( .A(decoded_rs2_2_bF_buf2_), .B(_6221_), .C(_6229_), .Y(_6230_) );
OAI21X1 OAI21X1_723 ( .A(_6215_), .B(decoded_rs2_3_bF_buf6_), .C(_6230_), .Y(_6231_) );
NOR2X1 NOR2X1_320 ( .A(_5347_), .B(_6231_), .Y(_6232_) );
NOR2X1 NOR2X1_321 ( .A(_5890__bF_buf2), .B(_6232_), .Y(_6233_) );
OAI21X1 OAI21X1_724 ( .A(decoded_rs2_4_bF_buf7_), .B(_6200_), .C(_6233_), .Y(_6234_) );
AOI21X1 AOI21X1_106 ( .A(decoded_imm_10_), .B(_5849__bF_buf4), .C(_4540__bF_buf2), .Y(_6235_) );
AOI22X1 AOI22X1_21 ( .A(_5122_), .B(_4540__bF_buf1), .C(_6234_), .D(_6235_), .Y(_82__10_) );
INVX1 INVX1_404 ( .A(cpuregs_2_[11]), .Y(_6236_) );
AOI21X1 AOI21X1_107 ( .A(decoded_rs2_1_bF_buf1_), .B(_6236_), .C(decoded_rs2_0_bF_buf52_), .Y(_6237_) );
OAI21X1 OAI21X1_725 ( .A(decoded_rs2_1_bF_buf0_), .B(cpuregs_0_[11]), .C(_6237_), .Y(_6238_) );
NOR2X1 NOR2X1_322 ( .A(decoded_rs2_1_bF_buf45_), .B(cpuregs_1_[11]), .Y(_6239_) );
OAI21X1 OAI21X1_726 ( .A(_5349__bF_buf1), .B(cpuregs_3_[11]), .C(decoded_rs2_0_bF_buf51_), .Y(_6240_) );
OAI21X1 OAI21X1_727 ( .A(_6239_), .B(_6240_), .C(_6238_), .Y(_6241_) );
NOR2X1 NOR2X1_323 ( .A(decoded_rs2_2_bF_buf1_), .B(_6241_), .Y(_6242_) );
AOI21X1 AOI21X1_108 ( .A(decoded_rs2_1_bF_buf44_), .B(_5289_), .C(decoded_rs2_0_bF_buf50_), .Y(_6243_) );
OAI21X1 OAI21X1_728 ( .A(decoded_rs2_1_bF_buf43_), .B(cpuregs_4_[11]), .C(_6243_), .Y(_6244_) );
NOR2X1 NOR2X1_324 ( .A(cpuregs_5_[11]), .B(decoded_rs2_1_bF_buf42_), .Y(_6245_) );
OAI21X1 OAI21X1_729 ( .A(_5349__bF_buf0), .B(cpuregs_7_[11]), .C(decoded_rs2_0_bF_buf49_), .Y(_6246_) );
OAI21X1 OAI21X1_730 ( .A(_6245_), .B(_6246_), .C(_6244_), .Y(_6247_) );
OAI21X1 OAI21X1_731 ( .A(_6247_), .B(_5358__bF_buf11), .C(_5348__bF_buf2), .Y(_6248_) );
INVX1 INVX1_405 ( .A(cpuregs_13_[11]), .Y(_6249_) );
AOI21X1 AOI21X1_109 ( .A(decoded_rs2_0_bF_buf48_), .B(_6249_), .C(decoded_rs2_1_bF_buf41_), .Y(_6250_) );
OAI21X1 OAI21X1_732 ( .A(decoded_rs2_0_bF_buf47_), .B(cpuregs_12_[11]), .C(_6250_), .Y(_6251_) );
NOR2X1 NOR2X1_325 ( .A(cpuregs_15_[11]), .B(_5362__bF_buf1), .Y(_6252_) );
OAI21X1 OAI21X1_733 ( .A(decoded_rs2_0_bF_buf46_), .B(cpuregs_14_[11]), .C(decoded_rs2_1_bF_buf40_), .Y(_6253_) );
OAI21X1 OAI21X1_734 ( .A(_6252_), .B(_6253_), .C(_6251_), .Y(_6254_) );
NOR2X1 NOR2X1_326 ( .A(_5358__bF_buf10), .B(_6254_), .Y(_6255_) );
INVX1 INVX1_406 ( .A(cpuregs_9_[11]), .Y(_6256_) );
AOI21X1 AOI21X1_110 ( .A(decoded_rs2_0_bF_buf45_), .B(_6256_), .C(decoded_rs2_1_bF_buf39_), .Y(_6257_) );
OAI21X1 OAI21X1_735 ( .A(cpuregs_8_[11]), .B(decoded_rs2_0_bF_buf44_), .C(_6257_), .Y(_6258_) );
NOR2X1 NOR2X1_327 ( .A(cpuregs_11_[11]), .B(_5362__bF_buf0), .Y(_6259_) );
OAI21X1 OAI21X1_736 ( .A(decoded_rs2_0_bF_buf43_), .B(cpuregs_10_[11]), .C(decoded_rs2_1_bF_buf38_), .Y(_6260_) );
OAI21X1 OAI21X1_737 ( .A(_6259_), .B(_6260_), .C(_6258_), .Y(_6261_) );
OAI21X1 OAI21X1_738 ( .A(_6261_), .B(decoded_rs2_2_bF_buf0_), .C(decoded_rs2_3_bF_buf5_), .Y(_6262_) );
OAI22X1 OAI22X1_37 ( .A(_6248_), .B(_6242_), .C(_6255_), .D(_6262_), .Y(_6263_) );
INVX1 INVX1_407 ( .A(cpuregs_26_[11]), .Y(_6264_) );
OAI21X1 OAI21X1_739 ( .A(_6264_), .B(decoded_rs2_0_bF_buf42_), .C(decoded_rs2_1_bF_buf37_), .Y(_6265_) );
AOI21X1 AOI21X1_111 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_27_[11]), .C(_6265_), .Y(_6266_) );
AND2X2 AND2X2_27 ( .A(decoded_rs2_0_bF_buf40_), .B(cpuregs_25_[11]), .Y(_6267_) );
INVX1 INVX1_408 ( .A(cpuregs_24_[11]), .Y(_6268_) );
OAI21X1 OAI21X1_740 ( .A(_6268_), .B(decoded_rs2_0_bF_buf39_), .C(_5349__bF_buf11), .Y(_6269_) );
OAI21X1 OAI21X1_741 ( .A(_6269_), .B(_6267_), .C(_5358__bF_buf9), .Y(_6270_) );
INVX1 INVX1_409 ( .A(cpuregs_28_[11]), .Y(_6271_) );
NAND2X1 NAND2X1_364 ( .A(decoded_rs2_0_bF_buf38_), .B(cpuregs_29_[11]), .Y(_6272_) );
OAI21X1 OAI21X1_742 ( .A(_6271_), .B(decoded_rs2_0_bF_buf37_), .C(_6272_), .Y(_6273_) );
INVX1 INVX1_410 ( .A(cpuregs_30_[11]), .Y(_6274_) );
NAND2X1 NAND2X1_365 ( .A(decoded_rs2_0_bF_buf36_), .B(cpuregs_31_[11]), .Y(_6275_) );
OAI21X1 OAI21X1_743 ( .A(_6274_), .B(decoded_rs2_0_bF_buf35_), .C(_6275_), .Y(_6276_) );
MUX2X1 MUX2X1_81 ( .A(_6276_), .B(_6273_), .S(decoded_rs2_1_bF_buf36_), .Y(_6277_) );
OAI22X1 OAI22X1_38 ( .A(_6270_), .B(_6266_), .C(_6277_), .D(_5358__bF_buf8), .Y(_6278_) );
INVX1 INVX1_411 ( .A(cpuregs_16_[11]), .Y(_6279_) );
NAND2X1 NAND2X1_366 ( .A(decoded_rs2_0_bF_buf34_), .B(cpuregs_17_[11]), .Y(_6280_) );
OAI21X1 OAI21X1_744 ( .A(_6279_), .B(decoded_rs2_0_bF_buf33_), .C(_6280_), .Y(_6281_) );
INVX1 INVX1_412 ( .A(cpuregs_19_[11]), .Y(_6282_) );
OAI21X1 OAI21X1_745 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_18_[11]), .C(decoded_rs2_1_bF_buf35_), .Y(_6283_) );
AOI21X1 AOI21X1_112 ( .A(decoded_rs2_0_bF_buf31_), .B(_6282_), .C(_6283_), .Y(_6284_) );
AOI21X1 AOI21X1_113 ( .A(_5349__bF_buf10), .B(_6281_), .C(_6284_), .Y(_6285_) );
NAND2X1 NAND2X1_367 ( .A(_5358__bF_buf7), .B(_6285_), .Y(_6286_) );
INVX1 INVX1_413 ( .A(cpuregs_20_[11]), .Y(_6287_) );
NAND2X1 NAND2X1_368 ( .A(decoded_rs2_0_bF_buf30_), .B(cpuregs_21_[11]), .Y(_6288_) );
OAI21X1 OAI21X1_746 ( .A(_6287_), .B(decoded_rs2_0_bF_buf29_), .C(_6288_), .Y(_6289_) );
INVX1 INVX1_414 ( .A(cpuregs_22_[11]), .Y(_6290_) );
NAND2X1 NAND2X1_369 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_23_[11]), .Y(_6291_) );
OAI21X1 OAI21X1_747 ( .A(_6290_), .B(decoded_rs2_0_bF_buf27_), .C(_6291_), .Y(_6292_) );
MUX2X1 MUX2X1_82 ( .A(_6292_), .B(_6289_), .S(decoded_rs2_1_bF_buf34_), .Y(_6293_) );
AOI21X1 AOI21X1_114 ( .A(decoded_rs2_2_bF_buf8_), .B(_6293_), .C(decoded_rs2_3_bF_buf4_), .Y(_6294_) );
AOI22X1 AOI22X1_22 ( .A(_6294_), .B(_6286_), .C(decoded_rs2_3_bF_buf3_), .D(_6278_), .Y(_6295_) );
AOI21X1 AOI21X1_115 ( .A(decoded_rs2_4_bF_buf6_), .B(_6295_), .C(_5890__bF_buf1), .Y(_6296_) );
OAI21X1 OAI21X1_748 ( .A(decoded_rs2_4_bF_buf5_), .B(_6263_), .C(_6296_), .Y(_6297_) );
AOI21X1 AOI21X1_116 ( .A(decoded_imm_11_), .B(_5849__bF_buf3), .C(_4540__bF_buf0), .Y(_6298_) );
AOI22X1 AOI22X1_23 ( .A(_5118_), .B(_4540__bF_buf6), .C(_6297_), .D(_6298_), .Y(_82__11_) );
NOR2X1 NOR2X1_328 ( .A(_10735__12_), .B(_4539__bF_buf3), .Y(_6299_) );
NOR2X1 NOR2X1_329 ( .A(cpuregs_8_[12]), .B(decoded_rs2_0_bF_buf26_), .Y(_6300_) );
OAI21X1 OAI21X1_749 ( .A(_5362__bF_buf14), .B(cpuregs_9_[12]), .C(_5349__bF_buf9), .Y(_6301_) );
NOR2X1 NOR2X1_330 ( .A(cpuregs_11_[12]), .B(_5362__bF_buf13), .Y(_6302_) );
OAI21X1 OAI21X1_750 ( .A(decoded_rs2_0_bF_buf25_), .B(cpuregs_10_[12]), .C(decoded_rs2_1_bF_buf33_), .Y(_6303_) );
OAI22X1 OAI22X1_39 ( .A(_6302_), .B(_6303_), .C(_6301_), .D(_6300_), .Y(_6304_) );
NOR2X1 NOR2X1_331 ( .A(decoded_rs2_0_bF_buf24_), .B(cpuregs_12_[12]), .Y(_6305_) );
OAI21X1 OAI21X1_751 ( .A(_5362__bF_buf12), .B(cpuregs_13_[12]), .C(_5349__bF_buf8), .Y(_6306_) );
NOR2X1 NOR2X1_332 ( .A(cpuregs_15_[12]), .B(_5362__bF_buf11), .Y(_6307_) );
OAI21X1 OAI21X1_752 ( .A(decoded_rs2_0_bF_buf23_), .B(cpuregs_14_[12]), .C(decoded_rs2_1_bF_buf32_), .Y(_6308_) );
OAI22X1 OAI22X1_40 ( .A(_6307_), .B(_6308_), .C(_6306_), .D(_6305_), .Y(_6309_) );
MUX2X1 MUX2X1_83 ( .A(_6309_), .B(_6304_), .S(decoded_rs2_2_bF_buf7_), .Y(_6310_) );
INVX1 INVX1_415 ( .A(cpuregs_6_[12]), .Y(_6311_) );
AOI21X1 AOI21X1_117 ( .A(decoded_rs2_1_bF_buf31_), .B(_6311_), .C(decoded_rs2_0_bF_buf22_), .Y(_6312_) );
OAI21X1 OAI21X1_753 ( .A(decoded_rs2_1_bF_buf30_), .B(cpuregs_4_[12]), .C(_6312_), .Y(_6313_) );
NOR2X1 NOR2X1_333 ( .A(cpuregs_5_[12]), .B(decoded_rs2_1_bF_buf29_), .Y(_6314_) );
OAI21X1 OAI21X1_754 ( .A(_5349__bF_buf7), .B(cpuregs_7_[12]), .C(decoded_rs2_0_bF_buf21_), .Y(_6315_) );
OAI21X1 OAI21X1_755 ( .A(_6314_), .B(_6315_), .C(_6313_), .Y(_6316_) );
INVX1 INVX1_416 ( .A(cpuregs_2_[12]), .Y(_6317_) );
AOI21X1 AOI21X1_118 ( .A(decoded_rs2_1_bF_buf28_), .B(_6317_), .C(decoded_rs2_0_bF_buf20_), .Y(_6318_) );
OAI21X1 OAI21X1_756 ( .A(decoded_rs2_1_bF_buf27_), .B(cpuregs_0_[12]), .C(_6318_), .Y(_6319_) );
NOR2X1 NOR2X1_334 ( .A(decoded_rs2_1_bF_buf26_), .B(cpuregs_1_[12]), .Y(_6320_) );
OAI21X1 OAI21X1_757 ( .A(_5349__bF_buf6), .B(cpuregs_3_[12]), .C(decoded_rs2_0_bF_buf19_), .Y(_6321_) );
OAI21X1 OAI21X1_758 ( .A(_6320_), .B(_6321_), .C(_6319_), .Y(_6322_) );
MUX2X1 MUX2X1_84 ( .A(_6322_), .B(_6316_), .S(_5358__bF_buf6), .Y(_6323_) );
MUX2X1 MUX2X1_85 ( .A(_6323_), .B(_6310_), .S(_5348__bF_buf1), .Y(_6324_) );
INVX1 INVX1_417 ( .A(cpuregs_16_[12]), .Y(_6325_) );
NAND2X1 NAND2X1_370 ( .A(decoded_rs2_0_bF_buf18_), .B(cpuregs_17_[12]), .Y(_6326_) );
OAI21X1 OAI21X1_759 ( .A(_6325_), .B(decoded_rs2_0_bF_buf17_), .C(_6326_), .Y(_6327_) );
INVX1 INVX1_418 ( .A(cpuregs_19_[12]), .Y(_6328_) );
OAI21X1 OAI21X1_760 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_18_[12]), .C(decoded_rs2_1_bF_buf25_), .Y(_6329_) );
AOI21X1 AOI21X1_119 ( .A(decoded_rs2_0_bF_buf15_), .B(_6328_), .C(_6329_), .Y(_6330_) );
AOI21X1 AOI21X1_120 ( .A(_5349__bF_buf5), .B(_6327_), .C(_6330_), .Y(_6331_) );
INVX1 INVX1_419 ( .A(cpuregs_20_[12]), .Y(_6332_) );
NAND2X1 NAND2X1_371 ( .A(decoded_rs2_0_bF_buf14_), .B(cpuregs_21_[12]), .Y(_6333_) );
OAI21X1 OAI21X1_761 ( .A(_6332_), .B(decoded_rs2_0_bF_buf13_), .C(_6333_), .Y(_6334_) );
INVX1 INVX1_420 ( .A(cpuregs_22_[12]), .Y(_6335_) );
NAND2X1 NAND2X1_372 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_23_[12]), .Y(_6336_) );
OAI21X1 OAI21X1_762 ( .A(_6335_), .B(decoded_rs2_0_bF_buf11_), .C(_6336_), .Y(_6337_) );
MUX2X1 MUX2X1_86 ( .A(_6337_), .B(_6334_), .S(decoded_rs2_1_bF_buf24_), .Y(_6338_) );
MUX2X1 MUX2X1_87 ( .A(_6331_), .B(_6338_), .S(_5358__bF_buf5), .Y(_6339_) );
NOR2X1 NOR2X1_335 ( .A(decoded_rs2_0_bF_buf10_), .B(cpuregs_24_[12]), .Y(_6340_) );
OAI21X1 OAI21X1_763 ( .A(_5362__bF_buf10), .B(cpuregs_25_[12]), .C(_5349__bF_buf4), .Y(_6341_) );
NOR2X1 NOR2X1_336 ( .A(_6340_), .B(_6341_), .Y(_6342_) );
INVX1 INVX1_421 ( .A(cpuregs_27_[12]), .Y(_6343_) );
OAI21X1 OAI21X1_764 ( .A(decoded_rs2_0_bF_buf9_), .B(cpuregs_26_[12]), .C(decoded_rs2_1_bF_buf23_), .Y(_6344_) );
AOI21X1 AOI21X1_121 ( .A(decoded_rs2_0_bF_buf8_), .B(_6343_), .C(_6344_), .Y(_6345_) );
OAI21X1 OAI21X1_765 ( .A(_6342_), .B(_6345_), .C(_5358__bF_buf4), .Y(_6346_) );
INVX1 INVX1_422 ( .A(cpuregs_28_[12]), .Y(_6347_) );
OAI21X1 OAI21X1_766 ( .A(_5362__bF_buf9), .B(cpuregs_29_[12]), .C(_5349__bF_buf3), .Y(_6348_) );
AOI21X1 AOI21X1_122 ( .A(_5362__bF_buf8), .B(_6347_), .C(_6348_), .Y(_6349_) );
INVX1 INVX1_423 ( .A(cpuregs_31_[12]), .Y(_6350_) );
OAI21X1 OAI21X1_767 ( .A(decoded_rs2_0_bF_buf7_), .B(cpuregs_30_[12]), .C(decoded_rs2_1_bF_buf22_), .Y(_6351_) );
AOI21X1 AOI21X1_123 ( .A(decoded_rs2_0_bF_buf6_), .B(_6350_), .C(_6351_), .Y(_6352_) );
OAI21X1 OAI21X1_768 ( .A(_6349_), .B(_6352_), .C(decoded_rs2_2_bF_buf6_), .Y(_6353_) );
AOI21X1 AOI21X1_124 ( .A(_6346_), .B(_6353_), .C(_5348__bF_buf0), .Y(_6354_) );
AOI21X1 AOI21X1_125 ( .A(_5348__bF_buf5), .B(_6339_), .C(_6354_), .Y(_6355_) );
AOI21X1 AOI21X1_126 ( .A(decoded_rs2_4_bF_buf4_), .B(_6355_), .C(_5890__bF_buf0), .Y(_6356_) );
OAI21X1 OAI21X1_769 ( .A(decoded_rs2_4_bF_buf3_), .B(_6324_), .C(_6356_), .Y(_6357_) );
AOI21X1 AOI21X1_127 ( .A(decoded_imm_12_), .B(_5849__bF_buf2), .C(_4540__bF_buf5), .Y(_6358_) );
AOI21X1 AOI21X1_128 ( .A(_6358_), .B(_6357_), .C(_6299_), .Y(_82__12_) );
NOR2X1 NOR2X1_337 ( .A(_10735__13_), .B(_4539__bF_buf2), .Y(_6359_) );
INVX1 INVX1_424 ( .A(cpuregs_9_[13]), .Y(_6360_) );
AOI21X1 AOI21X1_129 ( .A(decoded_rs2_0_bF_buf5_), .B(_6360_), .C(decoded_rs2_1_bF_buf21_), .Y(_6361_) );
OAI21X1 OAI21X1_770 ( .A(cpuregs_8_[13]), .B(decoded_rs2_0_bF_buf4_), .C(_6361_), .Y(_6362_) );
NOR2X1 NOR2X1_338 ( .A(cpuregs_11_[13]), .B(_5362__bF_buf7), .Y(_6363_) );
OAI21X1 OAI21X1_771 ( .A(decoded_rs2_0_bF_buf3_), .B(cpuregs_10_[13]), .C(decoded_rs2_1_bF_buf20_), .Y(_6364_) );
OAI21X1 OAI21X1_772 ( .A(_6363_), .B(_6364_), .C(_6362_), .Y(_6365_) );
INVX1 INVX1_425 ( .A(cpuregs_13_[13]), .Y(_6366_) );
AOI21X1 AOI21X1_130 ( .A(decoded_rs2_0_bF_buf2_), .B(_6366_), .C(decoded_rs2_1_bF_buf19_), .Y(_6367_) );
OAI21X1 OAI21X1_773 ( .A(decoded_rs2_0_bF_buf1_), .B(cpuregs_12_[13]), .C(_6367_), .Y(_6368_) );
NOR2X1 NOR2X1_339 ( .A(cpuregs_15_[13]), .B(_5362__bF_buf6), .Y(_6369_) );
OAI21X1 OAI21X1_774 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_14_[13]), .C(decoded_rs2_1_bF_buf18_), .Y(_6370_) );
OAI21X1 OAI21X1_775 ( .A(_6369_), .B(_6370_), .C(_6368_), .Y(_6371_) );
MUX2X1 MUX2X1_88 ( .A(_6371_), .B(_6365_), .S(decoded_rs2_2_bF_buf5_), .Y(_6372_) );
NOR2X1 NOR2X1_340 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_4_[13]), .Y(_6373_) );
OAI21X1 OAI21X1_776 ( .A(_5362__bF_buf5), .B(cpuregs_5_[13]), .C(_5349__bF_buf2), .Y(_6374_) );
NOR2X1 NOR2X1_341 ( .A(cpuregs_7_[13]), .B(_5362__bF_buf4), .Y(_6375_) );
OAI21X1 OAI21X1_777 ( .A(cpuregs_6_[13]), .B(decoded_rs2_0_bF_buf77_), .C(decoded_rs2_1_bF_buf17_), .Y(_6376_) );
OAI22X1 OAI22X1_41 ( .A(_6375_), .B(_6376_), .C(_6374_), .D(_6373_), .Y(_6377_) );
INVX1 INVX1_426 ( .A(cpuregs_2_[13]), .Y(_6378_) );
AOI21X1 AOI21X1_131 ( .A(decoded_rs2_1_bF_buf16_), .B(_6378_), .C(decoded_rs2_0_bF_buf76_), .Y(_6379_) );
OAI21X1 OAI21X1_778 ( .A(decoded_rs2_1_bF_buf15_), .B(cpuregs_0_[13]), .C(_6379_), .Y(_6380_) );
NOR2X1 NOR2X1_342 ( .A(decoded_rs2_1_bF_buf14_), .B(cpuregs_1_[13]), .Y(_6381_) );
OAI21X1 OAI21X1_779 ( .A(_5349__bF_buf1), .B(cpuregs_3_[13]), .C(decoded_rs2_0_bF_buf75_), .Y(_6382_) );
OAI21X1 OAI21X1_780 ( .A(_6381_), .B(_6382_), .C(_6380_), .Y(_6383_) );
MUX2X1 MUX2X1_89 ( .A(_6383_), .B(_6377_), .S(_5358__bF_buf3), .Y(_6384_) );
MUX2X1 MUX2X1_90 ( .A(_6372_), .B(_6384_), .S(decoded_rs2_3_bF_buf2_), .Y(_6385_) );
INVX1 INVX1_427 ( .A(cpuregs_16_[13]), .Y(_6386_) );
NAND2X1 NAND2X1_373 ( .A(decoded_rs2_0_bF_buf74_), .B(cpuregs_17_[13]), .Y(_6387_) );
OAI21X1 OAI21X1_781 ( .A(_6386_), .B(decoded_rs2_0_bF_buf73_), .C(_6387_), .Y(_6388_) );
INVX1 INVX1_428 ( .A(cpuregs_18_[13]), .Y(_6389_) );
NAND2X1 NAND2X1_374 ( .A(decoded_rs2_0_bF_buf72_), .B(cpuregs_19_[13]), .Y(_6390_) );
OAI21X1 OAI21X1_782 ( .A(_6389_), .B(decoded_rs2_0_bF_buf71_), .C(_6390_), .Y(_6391_) );
MUX2X1 MUX2X1_91 ( .A(_6391_), .B(_6388_), .S(decoded_rs2_1_bF_buf13_), .Y(_6392_) );
NOR2X1 NOR2X1_343 ( .A(decoded_rs2_2_bF_buf4_), .B(_6392_), .Y(_6393_) );
INVX1 INVX1_429 ( .A(cpuregs_20_[13]), .Y(_6394_) );
NAND2X1 NAND2X1_375 ( .A(decoded_rs2_0_bF_buf70_), .B(cpuregs_21_[13]), .Y(_6395_) );
OAI21X1 OAI21X1_783 ( .A(_6394_), .B(decoded_rs2_0_bF_buf69_), .C(_6395_), .Y(_6396_) );
INVX1 INVX1_430 ( .A(cpuregs_22_[13]), .Y(_6397_) );
NAND2X1 NAND2X1_376 ( .A(decoded_rs2_0_bF_buf68_), .B(cpuregs_23_[13]), .Y(_6398_) );
OAI21X1 OAI21X1_784 ( .A(_6397_), .B(decoded_rs2_0_bF_buf67_), .C(_6398_), .Y(_6399_) );
MUX2X1 MUX2X1_92 ( .A(_6399_), .B(_6396_), .S(decoded_rs2_1_bF_buf12_), .Y(_6400_) );
NOR2X1 NOR2X1_344 ( .A(_5358__bF_buf2), .B(_6400_), .Y(_6401_) );
OAI21X1 OAI21X1_785 ( .A(_6393_), .B(_6401_), .C(_5348__bF_buf4), .Y(_6402_) );
NOR2X1 NOR2X1_345 ( .A(decoded_rs2_0_bF_buf66_), .B(cpuregs_24_[13]), .Y(_6403_) );
OAI21X1 OAI21X1_786 ( .A(_5362__bF_buf3), .B(cpuregs_25_[13]), .C(_5349__bF_buf0), .Y(_6404_) );
NOR2X1 NOR2X1_346 ( .A(cpuregs_27_[13]), .B(_5362__bF_buf2), .Y(_6405_) );
OAI21X1 OAI21X1_787 ( .A(decoded_rs2_0_bF_buf65_), .B(cpuregs_26_[13]), .C(decoded_rs2_1_bF_buf11_), .Y(_6406_) );
OAI22X1 OAI22X1_42 ( .A(_6405_), .B(_6406_), .C(_6404_), .D(_6403_), .Y(_6407_) );
NOR2X1 NOR2X1_347 ( .A(decoded_rs2_2_bF_buf3_), .B(_6407_), .Y(_6408_) );
INVX1 INVX1_431 ( .A(cpuregs_29_[13]), .Y(_6409_) );
AOI21X1 AOI21X1_132 ( .A(decoded_rs2_0_bF_buf64_), .B(_6409_), .C(decoded_rs2_1_bF_buf10_), .Y(_6410_) );
OAI21X1 OAI21X1_788 ( .A(decoded_rs2_0_bF_buf63_), .B(cpuregs_28_[13]), .C(_6410_), .Y(_6411_) );
NOR2X1 NOR2X1_348 ( .A(cpuregs_31_[13]), .B(_5362__bF_buf1), .Y(_6412_) );
OAI21X1 OAI21X1_789 ( .A(decoded_rs2_0_bF_buf62_), .B(cpuregs_30_[13]), .C(decoded_rs2_1_bF_buf9_), .Y(_6413_) );
OAI21X1 OAI21X1_790 ( .A(_6412_), .B(_6413_), .C(_6411_), .Y(_6414_) );
OAI21X1 OAI21X1_791 ( .A(_6414_), .B(_5358__bF_buf1), .C(decoded_rs2_3_bF_buf1_), .Y(_6415_) );
OAI21X1 OAI21X1_792 ( .A(_6408_), .B(_6415_), .C(_6402_), .Y(_6416_) );
NOR2X1 NOR2X1_349 ( .A(_5347_), .B(_6416_), .Y(_6417_) );
NOR2X1 NOR2X1_350 ( .A(_5890__bF_buf3), .B(_6417_), .Y(_6418_) );
OAI21X1 OAI21X1_793 ( .A(decoded_rs2_4_bF_buf2_), .B(_6385_), .C(_6418_), .Y(_6419_) );
AOI21X1 AOI21X1_133 ( .A(decoded_imm_13_), .B(_5849__bF_buf1), .C(_4540__bF_buf4), .Y(_6420_) );
AOI21X1 AOI21X1_134 ( .A(_6420_), .B(_6419_), .C(_6359_), .Y(_82__13_) );
NOR2X1 NOR2X1_351 ( .A(_10735__14_), .B(_4539__bF_buf1), .Y(_6421_) );
INVX1 INVX1_432 ( .A(_5890__bF_buf2), .Y(_6422_) );
INVX1 INVX1_433 ( .A(cpuregs_20_[14]), .Y(_6423_) );
OAI21X1 OAI21X1_794 ( .A(_5358__bF_buf0), .B(_6423_), .C(_5362__bF_buf0), .Y(_6424_) );
AOI21X1 AOI21X1_135 ( .A(_5358__bF_buf12), .B(cpuregs_16_[14]), .C(_6424_), .Y(_6425_) );
INVX1 INVX1_434 ( .A(cpuregs_21_[14]), .Y(_6426_) );
OAI21X1 OAI21X1_795 ( .A(_5358__bF_buf11), .B(_6426_), .C(decoded_rs2_0_bF_buf61_), .Y(_6427_) );
AOI21X1 AOI21X1_136 ( .A(_5358__bF_buf10), .B(cpuregs_17_[14]), .C(_6427_), .Y(_6428_) );
OAI21X1 OAI21X1_796 ( .A(_6425_), .B(_6428_), .C(_5349__bF_buf11), .Y(_6429_) );
INVX1 INVX1_435 ( .A(cpuregs_22_[14]), .Y(_6430_) );
OAI21X1 OAI21X1_797 ( .A(_5358__bF_buf9), .B(_6430_), .C(_5362__bF_buf14), .Y(_6431_) );
AOI21X1 AOI21X1_137 ( .A(_5358__bF_buf8), .B(cpuregs_18_[14]), .C(_6431_), .Y(_6432_) );
INVX1 INVX1_436 ( .A(cpuregs_23_[14]), .Y(_6433_) );
OAI21X1 OAI21X1_798 ( .A(_5358__bF_buf7), .B(_6433_), .C(decoded_rs2_0_bF_buf60_), .Y(_6434_) );
AOI21X1 AOI21X1_138 ( .A(_5358__bF_buf6), .B(cpuregs_19_[14]), .C(_6434_), .Y(_6435_) );
OAI21X1 OAI21X1_799 ( .A(_6432_), .B(_6435_), .C(decoded_rs2_1_bF_buf8_), .Y(_6436_) );
NAND3X1 NAND3X1_22 ( .A(decoded_rs2_4_bF_buf1_), .B(_6429_), .C(_6436_), .Y(_6437_) );
NOR2X1 NOR2X1_352 ( .A(decoded_rs2_0_bF_buf59_), .B(cpuregs_4_[14]), .Y(_6438_) );
OAI21X1 OAI21X1_800 ( .A(_5362__bF_buf13), .B(cpuregs_5_[14]), .C(_5349__bF_buf10), .Y(_6439_) );
NOR2X1 NOR2X1_353 ( .A(cpuregs_7_[14]), .B(_5362__bF_buf12), .Y(_6440_) );
OAI21X1 OAI21X1_801 ( .A(cpuregs_6_[14]), .B(decoded_rs2_0_bF_buf58_), .C(decoded_rs2_1_bF_buf7_), .Y(_6441_) );
OAI22X1 OAI22X1_43 ( .A(_6440_), .B(_6441_), .C(_6439_), .D(_6438_), .Y(_6442_) );
NOR2X1 NOR2X1_354 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_0_[14]), .Y(_6443_) );
OAI21X1 OAI21X1_802 ( .A(_5362__bF_buf11), .B(cpuregs_1_[14]), .C(_5349__bF_buf9), .Y(_6444_) );
NOR2X1 NOR2X1_355 ( .A(cpuregs_3_[14]), .B(_5362__bF_buf10), .Y(_6445_) );
OAI21X1 OAI21X1_803 ( .A(decoded_rs2_0_bF_buf56_), .B(cpuregs_2_[14]), .C(decoded_rs2_1_bF_buf6_), .Y(_6446_) );
OAI22X1 OAI22X1_44 ( .A(_6445_), .B(_6446_), .C(_6444_), .D(_6443_), .Y(_6447_) );
MUX2X1 MUX2X1_93 ( .A(_6447_), .B(_6442_), .S(_5358__bF_buf5), .Y(_6448_) );
OAI21X1 OAI21X1_804 ( .A(decoded_rs2_4_bF_buf0_), .B(_6448_), .C(_6437_), .Y(_6449_) );
AND2X2 AND2X2_28 ( .A(_6449_), .B(_5348__bF_buf3), .Y(_6450_) );
INVX1 INVX1_437 ( .A(cpuregs_28_[14]), .Y(_6451_) );
NAND2X1 NAND2X1_377 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_29_[14]), .Y(_6452_) );
OAI21X1 OAI21X1_805 ( .A(_6451_), .B(decoded_rs2_0_bF_buf54_), .C(_6452_), .Y(_6453_) );
INVX1 INVX1_438 ( .A(cpuregs_31_[14]), .Y(_6454_) );
OAI21X1 OAI21X1_806 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_30_[14]), .C(decoded_rs2_1_bF_buf5_), .Y(_6455_) );
AOI21X1 AOI21X1_139 ( .A(decoded_rs2_0_bF_buf52_), .B(_6454_), .C(_6455_), .Y(_6456_) );
AOI21X1 AOI21X1_140 ( .A(_5349__bF_buf8), .B(_6453_), .C(_6456_), .Y(_6457_) );
NOR2X1 NOR2X1_356 ( .A(_5358__bF_buf4), .B(_6457_), .Y(_6458_) );
INVX1 INVX1_439 ( .A(cpuregs_24_[14]), .Y(_6459_) );
NAND2X1 NAND2X1_378 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_25_[14]), .Y(_6460_) );
OAI21X1 OAI21X1_807 ( .A(_6459_), .B(decoded_rs2_0_bF_buf50_), .C(_6460_), .Y(_6461_) );
INVX1 INVX1_440 ( .A(cpuregs_27_[14]), .Y(_6462_) );
OAI21X1 OAI21X1_808 ( .A(decoded_rs2_0_bF_buf49_), .B(cpuregs_26_[14]), .C(decoded_rs2_1_bF_buf4_), .Y(_6463_) );
AOI21X1 AOI21X1_141 ( .A(decoded_rs2_0_bF_buf48_), .B(_6462_), .C(_6463_), .Y(_6464_) );
AOI21X1 AOI21X1_142 ( .A(_5349__bF_buf7), .B(_6461_), .C(_6464_), .Y(_6465_) );
NOR2X1 NOR2X1_357 ( .A(decoded_rs2_2_bF_buf2_), .B(_6465_), .Y(_6466_) );
OAI21X1 OAI21X1_809 ( .A(_6458_), .B(_6466_), .C(decoded_rs2_4_bF_buf7_), .Y(_6467_) );
INVX1 INVX1_441 ( .A(cpuregs_9_[14]), .Y(_6468_) );
AOI21X1 AOI21X1_143 ( .A(decoded_rs2_0_bF_buf47_), .B(_6468_), .C(decoded_rs2_1_bF_buf3_), .Y(_6469_) );
OAI21X1 OAI21X1_810 ( .A(cpuregs_8_[14]), .B(decoded_rs2_0_bF_buf46_), .C(_6469_), .Y(_6470_) );
NOR2X1 NOR2X1_358 ( .A(cpuregs_11_[14]), .B(_5362__bF_buf9), .Y(_6471_) );
OAI21X1 OAI21X1_811 ( .A(decoded_rs2_0_bF_buf45_), .B(cpuregs_10_[14]), .C(decoded_rs2_1_bF_buf2_), .Y(_6472_) );
OAI21X1 OAI21X1_812 ( .A(_6471_), .B(_6472_), .C(_6470_), .Y(_6473_) );
INVX1 INVX1_442 ( .A(cpuregs_13_[14]), .Y(_6474_) );
AOI21X1 AOI21X1_144 ( .A(decoded_rs2_0_bF_buf44_), .B(_6474_), .C(decoded_rs2_1_bF_buf1_), .Y(_6475_) );
OAI21X1 OAI21X1_813 ( .A(decoded_rs2_0_bF_buf43_), .B(cpuregs_12_[14]), .C(_6475_), .Y(_6476_) );
NOR2X1 NOR2X1_359 ( .A(cpuregs_15_[14]), .B(_5362__bF_buf8), .Y(_6477_) );
OAI21X1 OAI21X1_814 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_14_[14]), .C(decoded_rs2_1_bF_buf0_), .Y(_6478_) );
OAI21X1 OAI21X1_815 ( .A(_6477_), .B(_6478_), .C(_6476_), .Y(_6479_) );
MUX2X1 MUX2X1_94 ( .A(_6479_), .B(_6473_), .S(decoded_rs2_2_bF_buf1_), .Y(_6480_) );
OAI21X1 OAI21X1_816 ( .A(decoded_rs2_4_bF_buf6_), .B(_6480_), .C(_6467_), .Y(_6481_) );
AND2X2 AND2X2_29 ( .A(_6481_), .B(decoded_rs2_3_bF_buf0_), .Y(_6482_) );
OAI21X1 OAI21X1_817 ( .A(_6482_), .B(_6450_), .C(_6422_), .Y(_6483_) );
AOI21X1 AOI21X1_145 ( .A(decoded_imm_14_), .B(_5849__bF_buf0), .C(_4540__bF_buf3), .Y(_6484_) );
AOI21X1 AOI21X1_146 ( .A(_6484_), .B(_6483_), .C(_6421_), .Y(_82__14_) );
NOR2X1 NOR2X1_360 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_4_[15]), .Y(_6485_) );
OAI21X1 OAI21X1_818 ( .A(_5362__bF_buf7), .B(cpuregs_5_[15]), .C(_5349__bF_buf6), .Y(_6486_) );
NOR2X1 NOR2X1_361 ( .A(cpuregs_7_[15]), .B(_5362__bF_buf6), .Y(_6487_) );
OAI21X1 OAI21X1_819 ( .A(cpuregs_6_[15]), .B(decoded_rs2_0_bF_buf40_), .C(decoded_rs2_1_bF_buf45_), .Y(_6488_) );
OAI22X1 OAI22X1_45 ( .A(_6487_), .B(_6488_), .C(_6486_), .D(_6485_), .Y(_6489_) );
INVX1 INVX1_443 ( .A(cpuregs_2_[15]), .Y(_6490_) );
AOI21X1 AOI21X1_147 ( .A(decoded_rs2_1_bF_buf44_), .B(_6490_), .C(decoded_rs2_0_bF_buf39_), .Y(_6491_) );
OAI21X1 OAI21X1_820 ( .A(decoded_rs2_1_bF_buf43_), .B(cpuregs_0_[15]), .C(_6491_), .Y(_6492_) );
NOR2X1 NOR2X1_362 ( .A(decoded_rs2_1_bF_buf42_), .B(cpuregs_1_[15]), .Y(_6493_) );
OAI21X1 OAI21X1_821 ( .A(_5349__bF_buf5), .B(cpuregs_3_[15]), .C(decoded_rs2_0_bF_buf38_), .Y(_6494_) );
OAI21X1 OAI21X1_822 ( .A(_6493_), .B(_6494_), .C(_6492_), .Y(_6495_) );
MUX2X1 MUX2X1_95 ( .A(_6495_), .B(_6489_), .S(_5358__bF_buf3), .Y(_6496_) );
INVX1 INVX1_444 ( .A(cpuregs_9_[15]), .Y(_6497_) );
AOI21X1 AOI21X1_148 ( .A(decoded_rs2_0_bF_buf37_), .B(_6497_), .C(decoded_rs2_1_bF_buf41_), .Y(_6498_) );
OAI21X1 OAI21X1_823 ( .A(cpuregs_8_[15]), .B(decoded_rs2_0_bF_buf36_), .C(_6498_), .Y(_6499_) );
NOR2X1 NOR2X1_363 ( .A(cpuregs_11_[15]), .B(_5362__bF_buf5), .Y(_6500_) );
OAI21X1 OAI21X1_824 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_10_[15]), .C(decoded_rs2_1_bF_buf40_), .Y(_6501_) );
OAI21X1 OAI21X1_825 ( .A(_6500_), .B(_6501_), .C(_6499_), .Y(_6502_) );
INVX1 INVX1_445 ( .A(cpuregs_13_[15]), .Y(_6503_) );
AOI21X1 AOI21X1_149 ( .A(decoded_rs2_0_bF_buf34_), .B(_6503_), .C(decoded_rs2_1_bF_buf39_), .Y(_6504_) );
OAI21X1 OAI21X1_826 ( .A(decoded_rs2_0_bF_buf33_), .B(cpuregs_12_[15]), .C(_6504_), .Y(_6505_) );
NOR2X1 NOR2X1_364 ( .A(cpuregs_15_[15]), .B(_5362__bF_buf4), .Y(_6506_) );
OAI21X1 OAI21X1_827 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_14_[15]), .C(decoded_rs2_1_bF_buf38_), .Y(_6507_) );
OAI21X1 OAI21X1_828 ( .A(_6506_), .B(_6507_), .C(_6505_), .Y(_6508_) );
MUX2X1 MUX2X1_96 ( .A(_6508_), .B(_6502_), .S(decoded_rs2_2_bF_buf0_), .Y(_6509_) );
MUX2X1 MUX2X1_97 ( .A(_6509_), .B(_6496_), .S(decoded_rs2_3_bF_buf6_), .Y(_6510_) );
INVX1 INVX1_446 ( .A(cpuregs_28_[15]), .Y(_6511_) );
NAND2X1 NAND2X1_379 ( .A(decoded_rs2_0_bF_buf31_), .B(cpuregs_29_[15]), .Y(_6512_) );
OAI21X1 OAI21X1_829 ( .A(_6511_), .B(decoded_rs2_0_bF_buf30_), .C(_6512_), .Y(_6513_) );
INVX1 INVX1_447 ( .A(cpuregs_31_[15]), .Y(_6514_) );
OAI21X1 OAI21X1_830 ( .A(decoded_rs2_0_bF_buf29_), .B(cpuregs_30_[15]), .C(decoded_rs2_1_bF_buf37_), .Y(_6515_) );
AOI21X1 AOI21X1_150 ( .A(decoded_rs2_0_bF_buf28_), .B(_6514_), .C(_6515_), .Y(_6516_) );
AOI21X1 AOI21X1_151 ( .A(_5349__bF_buf4), .B(_6513_), .C(_6516_), .Y(_6517_) );
NOR2X1 NOR2X1_365 ( .A(_5358__bF_buf2), .B(_6517_), .Y(_6518_) );
INVX1 INVX1_448 ( .A(cpuregs_24_[15]), .Y(_6519_) );
NAND2X1 NAND2X1_380 ( .A(decoded_rs2_0_bF_buf27_), .B(cpuregs_25_[15]), .Y(_6520_) );
OAI21X1 OAI21X1_831 ( .A(_6519_), .B(decoded_rs2_0_bF_buf26_), .C(_6520_), .Y(_6521_) );
INVX1 INVX1_449 ( .A(cpuregs_27_[15]), .Y(_6522_) );
OAI21X1 OAI21X1_832 ( .A(decoded_rs2_0_bF_buf25_), .B(cpuregs_26_[15]), .C(decoded_rs2_1_bF_buf36_), .Y(_6523_) );
AOI21X1 AOI21X1_152 ( .A(decoded_rs2_0_bF_buf24_), .B(_6522_), .C(_6523_), .Y(_6524_) );
AOI21X1 AOI21X1_153 ( .A(_5349__bF_buf3), .B(_6521_), .C(_6524_), .Y(_6525_) );
NOR2X1 NOR2X1_366 ( .A(decoded_rs2_2_bF_buf8_), .B(_6525_), .Y(_6526_) );
OAI21X1 OAI21X1_833 ( .A(_6518_), .B(_6526_), .C(decoded_rs2_3_bF_buf5_), .Y(_6527_) );
INVX1 INVX1_450 ( .A(cpuregs_17_[15]), .Y(_6528_) );
AOI21X1 AOI21X1_154 ( .A(decoded_rs2_0_bF_buf23_), .B(_6528_), .C(decoded_rs2_1_bF_buf35_), .Y(_6529_) );
OAI21X1 OAI21X1_834 ( .A(decoded_rs2_0_bF_buf22_), .B(cpuregs_16_[15]), .C(_6529_), .Y(_6530_) );
NOR2X1 NOR2X1_367 ( .A(cpuregs_19_[15]), .B(_5362__bF_buf3), .Y(_6531_) );
OAI21X1 OAI21X1_835 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_18_[15]), .C(decoded_rs2_1_bF_buf34_), .Y(_6532_) );
OAI21X1 OAI21X1_836 ( .A(_6531_), .B(_6532_), .C(_6530_), .Y(_6533_) );
INVX1 INVX1_451 ( .A(cpuregs_21_[15]), .Y(_6534_) );
AOI21X1 AOI21X1_155 ( .A(decoded_rs2_0_bF_buf20_), .B(_6534_), .C(decoded_rs2_1_bF_buf33_), .Y(_6535_) );
OAI21X1 OAI21X1_837 ( .A(decoded_rs2_0_bF_buf19_), .B(cpuregs_20_[15]), .C(_6535_), .Y(_6536_) );
INVX1 INVX1_452 ( .A(cpuregs_22_[15]), .Y(_6537_) );
AOI21X1 AOI21X1_156 ( .A(_5362__bF_buf2), .B(_6537_), .C(_5349__bF_buf2), .Y(_6538_) );
OAI21X1 OAI21X1_838 ( .A(_5362__bF_buf1), .B(cpuregs_23_[15]), .C(_6538_), .Y(_6539_) );
NAND3X1 NAND3X1_23 ( .A(decoded_rs2_2_bF_buf7_), .B(_6536_), .C(_6539_), .Y(_6540_) );
OAI21X1 OAI21X1_839 ( .A(_6533_), .B(decoded_rs2_2_bF_buf6_), .C(_6540_), .Y(_6541_) );
OAI21X1 OAI21X1_840 ( .A(decoded_rs2_3_bF_buf4_), .B(_6541_), .C(_6527_), .Y(_6542_) );
NOR2X1 NOR2X1_368 ( .A(_5347_), .B(_6542_), .Y(_6543_) );
NOR2X1 NOR2X1_369 ( .A(_5890__bF_buf1), .B(_6543_), .Y(_6544_) );
OAI21X1 OAI21X1_841 ( .A(decoded_rs2_4_bF_buf5_), .B(_6510_), .C(_6544_), .Y(_6545_) );
AOI21X1 AOI21X1_157 ( .A(decoded_imm_15_), .B(_5849__bF_buf4), .C(_4540__bF_buf2), .Y(_6546_) );
AOI22X1 AOI22X1_24 ( .A(_5088_), .B(_4540__bF_buf1), .C(_6545_), .D(_6546_), .Y(_82__15_) );
INVX1 INVX1_453 ( .A(cpuregs_20_[16]), .Y(_6547_) );
OAI21X1 OAI21X1_842 ( .A(_5358__bF_buf1), .B(_6547_), .C(_5362__bF_buf0), .Y(_6548_) );
AOI21X1 AOI21X1_158 ( .A(_5358__bF_buf0), .B(cpuregs_16_[16]), .C(_6548_), .Y(_6549_) );
INVX1 INVX1_454 ( .A(cpuregs_21_[16]), .Y(_6550_) );
OAI21X1 OAI21X1_843 ( .A(_5358__bF_buf12), .B(_6550_), .C(decoded_rs2_0_bF_buf18_), .Y(_6551_) );
AOI21X1 AOI21X1_159 ( .A(_5358__bF_buf11), .B(cpuregs_17_[16]), .C(_6551_), .Y(_6552_) );
OAI21X1 OAI21X1_844 ( .A(_6549_), .B(_6552_), .C(_5349__bF_buf1), .Y(_6553_) );
INVX1 INVX1_455 ( .A(cpuregs_22_[16]), .Y(_6554_) );
OAI21X1 OAI21X1_845 ( .A(_5358__bF_buf10), .B(_6554_), .C(_5362__bF_buf14), .Y(_6555_) );
AOI21X1 AOI21X1_160 ( .A(_5358__bF_buf9), .B(cpuregs_18_[16]), .C(_6555_), .Y(_6556_) );
INVX1 INVX1_456 ( .A(cpuregs_23_[16]), .Y(_6557_) );
OAI21X1 OAI21X1_846 ( .A(_5358__bF_buf8), .B(_6557_), .C(decoded_rs2_0_bF_buf17_), .Y(_6558_) );
AOI21X1 AOI21X1_161 ( .A(_5358__bF_buf7), .B(cpuregs_19_[16]), .C(_6558_), .Y(_6559_) );
OAI21X1 OAI21X1_847 ( .A(_6556_), .B(_6559_), .C(decoded_rs2_1_bF_buf32_), .Y(_6560_) );
NAND3X1 NAND3X1_24 ( .A(decoded_rs2_4_bF_buf4_), .B(_6553_), .C(_6560_), .Y(_6561_) );
NOR2X1 NOR2X1_370 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_4_[16]), .Y(_6562_) );
OAI21X1 OAI21X1_848 ( .A(_5362__bF_buf13), .B(cpuregs_5_[16]), .C(_5349__bF_buf0), .Y(_6563_) );
NOR2X1 NOR2X1_371 ( .A(cpuregs_7_[16]), .B(_5362__bF_buf12), .Y(_6564_) );
OAI21X1 OAI21X1_849 ( .A(cpuregs_6_[16]), .B(decoded_rs2_0_bF_buf15_), .C(decoded_rs2_1_bF_buf31_), .Y(_6565_) );
OAI22X1 OAI22X1_46 ( .A(_6564_), .B(_6565_), .C(_6563_), .D(_6562_), .Y(_6566_) );
NOR2X1 NOR2X1_372 ( .A(decoded_rs2_0_bF_buf14_), .B(cpuregs_0_[16]), .Y(_6567_) );
OAI21X1 OAI21X1_850 ( .A(_5362__bF_buf11), .B(cpuregs_1_[16]), .C(_5349__bF_buf11), .Y(_6568_) );
NOR2X1 NOR2X1_373 ( .A(cpuregs_3_[16]), .B(_5362__bF_buf10), .Y(_6569_) );
OAI21X1 OAI21X1_851 ( .A(decoded_rs2_0_bF_buf13_), .B(cpuregs_2_[16]), .C(decoded_rs2_1_bF_buf30_), .Y(_6570_) );
OAI22X1 OAI22X1_47 ( .A(_6569_), .B(_6570_), .C(_6568_), .D(_6567_), .Y(_6571_) );
MUX2X1 MUX2X1_98 ( .A(_6571_), .B(_6566_), .S(_5358__bF_buf6), .Y(_6572_) );
OAI21X1 OAI21X1_852 ( .A(decoded_rs2_4_bF_buf3_), .B(_6572_), .C(_6561_), .Y(_6573_) );
AND2X2 AND2X2_30 ( .A(_6573_), .B(_5348__bF_buf2), .Y(_6574_) );
INVX1 INVX1_457 ( .A(cpuregs_29_[16]), .Y(_6575_) );
NAND2X1 NAND2X1_381 ( .A(cpuregs_28_[16]), .B(_5362__bF_buf9), .Y(_6576_) );
OAI21X1 OAI21X1_853 ( .A(_5362__bF_buf8), .B(_6575_), .C(_6576_), .Y(_6577_) );
INVX1 INVX1_458 ( .A(cpuregs_31_[16]), .Y(_6578_) );
OAI21X1 OAI21X1_854 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_30_[16]), .C(decoded_rs2_1_bF_buf29_), .Y(_6579_) );
AOI21X1 AOI21X1_162 ( .A(decoded_rs2_0_bF_buf11_), .B(_6578_), .C(_6579_), .Y(_6580_) );
AOI21X1 AOI21X1_163 ( .A(_5349__bF_buf10), .B(_6577_), .C(_6580_), .Y(_6581_) );
NOR2X1 NOR2X1_374 ( .A(_5358__bF_buf5), .B(_6581_), .Y(_6582_) );
INVX1 INVX1_459 ( .A(cpuregs_24_[16]), .Y(_6583_) );
NAND2X1 NAND2X1_382 ( .A(decoded_rs2_0_bF_buf10_), .B(cpuregs_25_[16]), .Y(_6584_) );
OAI21X1 OAI21X1_855 ( .A(_6583_), .B(decoded_rs2_0_bF_buf9_), .C(_6584_), .Y(_6585_) );
INVX1 INVX1_460 ( .A(cpuregs_27_[16]), .Y(_6586_) );
OAI21X1 OAI21X1_856 ( .A(decoded_rs2_0_bF_buf8_), .B(cpuregs_26_[16]), .C(decoded_rs2_1_bF_buf28_), .Y(_6587_) );
AOI21X1 AOI21X1_164 ( .A(decoded_rs2_0_bF_buf7_), .B(_6586_), .C(_6587_), .Y(_6588_) );
AOI21X1 AOI21X1_165 ( .A(_5349__bF_buf9), .B(_6585_), .C(_6588_), .Y(_6589_) );
NOR2X1 NOR2X1_375 ( .A(decoded_rs2_2_bF_buf5_), .B(_6589_), .Y(_6590_) );
OAI21X1 OAI21X1_857 ( .A(_6582_), .B(_6590_), .C(decoded_rs2_4_bF_buf2_), .Y(_6591_) );
NOR2X1 NOR2X1_376 ( .A(cpuregs_8_[16]), .B(decoded_rs2_0_bF_buf6_), .Y(_6592_) );
OAI21X1 OAI21X1_858 ( .A(_5362__bF_buf7), .B(cpuregs_9_[16]), .C(_5349__bF_buf8), .Y(_6593_) );
NOR2X1 NOR2X1_377 ( .A(cpuregs_11_[16]), .B(_5362__bF_buf6), .Y(_6594_) );
OAI21X1 OAI21X1_859 ( .A(decoded_rs2_0_bF_buf5_), .B(cpuregs_10_[16]), .C(decoded_rs2_1_bF_buf27_), .Y(_6595_) );
OAI22X1 OAI22X1_48 ( .A(_6594_), .B(_6595_), .C(_6593_), .D(_6592_), .Y(_6596_) );
NOR2X1 NOR2X1_378 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_12_[16]), .Y(_6597_) );
OAI21X1 OAI21X1_860 ( .A(_5362__bF_buf5), .B(cpuregs_13_[16]), .C(_5349__bF_buf7), .Y(_6598_) );
NOR2X1 NOR2X1_379 ( .A(cpuregs_15_[16]), .B(_5362__bF_buf4), .Y(_6599_) );
OAI21X1 OAI21X1_861 ( .A(decoded_rs2_0_bF_buf3_), .B(cpuregs_14_[16]), .C(decoded_rs2_1_bF_buf26_), .Y(_6600_) );
OAI22X1 OAI22X1_49 ( .A(_6599_), .B(_6600_), .C(_6598_), .D(_6597_), .Y(_6601_) );
MUX2X1 MUX2X1_99 ( .A(_6596_), .B(_6601_), .S(_5358__bF_buf4), .Y(_6602_) );
OAI21X1 OAI21X1_862 ( .A(decoded_rs2_4_bF_buf1_), .B(_6602_), .C(_6591_), .Y(_6603_) );
AND2X2 AND2X2_31 ( .A(_6603_), .B(decoded_rs2_3_bF_buf3_), .Y(_6604_) );
OAI21X1 OAI21X1_863 ( .A(_6604_), .B(_6574_), .C(_6422_), .Y(_6605_) );
AOI21X1 AOI21X1_166 ( .A(decoded_imm_16_), .B(_5849__bF_buf3), .C(_4540__bF_buf0), .Y(_6606_) );
AOI22X1 AOI22X1_25 ( .A(_5052_), .B(_4540__bF_buf6), .C(_6605_), .D(_6606_), .Y(_82__16_) );
INVX1 INVX1_461 ( .A(cpuregs_20_[17]), .Y(_6607_) );
OAI21X1 OAI21X1_864 ( .A(_5358__bF_buf3), .B(_6607_), .C(_5362__bF_buf3), .Y(_6608_) );
AOI21X1 AOI21X1_167 ( .A(_5358__bF_buf2), .B(cpuregs_16_[17]), .C(_6608_), .Y(_6609_) );
INVX1 INVX1_462 ( .A(cpuregs_21_[17]), .Y(_6610_) );
OAI21X1 OAI21X1_865 ( .A(_5358__bF_buf1), .B(_6610_), .C(decoded_rs2_0_bF_buf2_), .Y(_6611_) );
AOI21X1 AOI21X1_168 ( .A(_5358__bF_buf0), .B(cpuregs_17_[17]), .C(_6611_), .Y(_6612_) );
OAI21X1 OAI21X1_866 ( .A(_6609_), .B(_6612_), .C(_5349__bF_buf6), .Y(_6613_) );
INVX1 INVX1_463 ( .A(cpuregs_22_[17]), .Y(_6614_) );
OAI21X1 OAI21X1_867 ( .A(_5358__bF_buf12), .B(_6614_), .C(_5362__bF_buf2), .Y(_6615_) );
AOI21X1 AOI21X1_169 ( .A(_5358__bF_buf11), .B(cpuregs_18_[17]), .C(_6615_), .Y(_6616_) );
INVX1 INVX1_464 ( .A(cpuregs_23_[17]), .Y(_6617_) );
OAI21X1 OAI21X1_868 ( .A(_5358__bF_buf10), .B(_6617_), .C(decoded_rs2_0_bF_buf1_), .Y(_6618_) );
AOI21X1 AOI21X1_170 ( .A(_5358__bF_buf9), .B(cpuregs_19_[17]), .C(_6618_), .Y(_6619_) );
OAI21X1 OAI21X1_869 ( .A(_6616_), .B(_6619_), .C(decoded_rs2_1_bF_buf25_), .Y(_6620_) );
NAND3X1 NAND3X1_25 ( .A(decoded_rs2_4_bF_buf0_), .B(_6613_), .C(_6620_), .Y(_6621_) );
INVX1 INVX1_465 ( .A(cpuregs_0_[17]), .Y(_6622_) );
NAND2X1 NAND2X1_383 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_1_[17]), .Y(_6623_) );
OAI21X1 OAI21X1_870 ( .A(_6622_), .B(decoded_rs2_0_bF_buf78_), .C(_6623_), .Y(_6624_) );
INVX1 INVX1_466 ( .A(cpuregs_2_[17]), .Y(_6625_) );
NAND2X1 NAND2X1_384 ( .A(decoded_rs2_0_bF_buf77_), .B(cpuregs_3_[17]), .Y(_6626_) );
OAI21X1 OAI21X1_871 ( .A(_6625_), .B(decoded_rs2_0_bF_buf76_), .C(_6626_), .Y(_6627_) );
MUX2X1 MUX2X1_100 ( .A(_6627_), .B(_6624_), .S(decoded_rs2_1_bF_buf24_), .Y(_6628_) );
NAND2X1 NAND2X1_385 ( .A(_5358__bF_buf8), .B(_6628_), .Y(_6629_) );
NOR2X1 NOR2X1_380 ( .A(decoded_rs2_0_bF_buf75_), .B(cpuregs_4_[17]), .Y(_6630_) );
OAI21X1 OAI21X1_872 ( .A(_5362__bF_buf1), .B(cpuregs_5_[17]), .C(_5349__bF_buf5), .Y(_6631_) );
NOR2X1 NOR2X1_381 ( .A(cpuregs_7_[17]), .B(_5362__bF_buf0), .Y(_6632_) );
OAI21X1 OAI21X1_873 ( .A(cpuregs_6_[17]), .B(decoded_rs2_0_bF_buf74_), .C(decoded_rs2_1_bF_buf23_), .Y(_6633_) );
OAI22X1 OAI22X1_50 ( .A(_6632_), .B(_6633_), .C(_6631_), .D(_6630_), .Y(_6634_) );
OAI21X1 OAI21X1_874 ( .A(_5358__bF_buf7), .B(_6634_), .C(_6629_), .Y(_6635_) );
OAI21X1 OAI21X1_875 ( .A(decoded_rs2_4_bF_buf7_), .B(_6635_), .C(_6621_), .Y(_6636_) );
AND2X2 AND2X2_32 ( .A(_6636_), .B(_5348__bF_buf1), .Y(_6637_) );
INVX1 INVX1_467 ( .A(cpuregs_28_[17]), .Y(_6638_) );
NAND2X1 NAND2X1_386 ( .A(decoded_rs2_0_bF_buf73_), .B(cpuregs_29_[17]), .Y(_6639_) );
OAI21X1 OAI21X1_876 ( .A(_6638_), .B(decoded_rs2_0_bF_buf72_), .C(_6639_), .Y(_6640_) );
INVX1 INVX1_468 ( .A(cpuregs_31_[17]), .Y(_6641_) );
OAI21X1 OAI21X1_877 ( .A(decoded_rs2_0_bF_buf71_), .B(cpuregs_30_[17]), .C(decoded_rs2_1_bF_buf22_), .Y(_6642_) );
AOI21X1 AOI21X1_171 ( .A(decoded_rs2_0_bF_buf70_), .B(_6641_), .C(_6642_), .Y(_6643_) );
AOI21X1 AOI21X1_172 ( .A(_5349__bF_buf4), .B(_6640_), .C(_6643_), .Y(_6644_) );
INVX1 INVX1_469 ( .A(cpuregs_24_[17]), .Y(_6645_) );
NAND2X1 NAND2X1_387 ( .A(decoded_rs2_0_bF_buf69_), .B(cpuregs_25_[17]), .Y(_6646_) );
OAI21X1 OAI21X1_878 ( .A(_6645_), .B(decoded_rs2_0_bF_buf68_), .C(_6646_), .Y(_6647_) );
INVX1 INVX1_470 ( .A(cpuregs_27_[17]), .Y(_6648_) );
OAI21X1 OAI21X1_879 ( .A(decoded_rs2_0_bF_buf67_), .B(cpuregs_26_[17]), .C(decoded_rs2_1_bF_buf21_), .Y(_6649_) );
AOI21X1 AOI21X1_173 ( .A(decoded_rs2_0_bF_buf66_), .B(_6648_), .C(_6649_), .Y(_6650_) );
AOI21X1 AOI21X1_174 ( .A(_5349__bF_buf3), .B(_6647_), .C(_6650_), .Y(_6651_) );
MUX2X1 MUX2X1_101 ( .A(_6651_), .B(_6644_), .S(_5358__bF_buf6), .Y(_6652_) );
INVX1 INVX1_471 ( .A(cpuregs_9_[17]), .Y(_6653_) );
OAI21X1 OAI21X1_880 ( .A(_6653_), .B(decoded_rs2_1_bF_buf20_), .C(decoded_rs2_0_bF_buf65_), .Y(_6654_) );
AOI21X1 AOI21X1_175 ( .A(decoded_rs2_1_bF_buf19_), .B(cpuregs_11_[17]), .C(_6654_), .Y(_6655_) );
AND2X2 AND2X2_33 ( .A(decoded_rs2_1_bF_buf18_), .B(cpuregs_10_[17]), .Y(_6656_) );
INVX1 INVX1_472 ( .A(cpuregs_8_[17]), .Y(_6657_) );
OAI21X1 OAI21X1_881 ( .A(_6657_), .B(decoded_rs2_1_bF_buf17_), .C(_5362__bF_buf14), .Y(_6658_) );
OAI21X1 OAI21X1_882 ( .A(_6658_), .B(_6656_), .C(_5358__bF_buf5), .Y(_6659_) );
INVX1 INVX1_473 ( .A(cpuregs_13_[17]), .Y(_6660_) );
OAI21X1 OAI21X1_883 ( .A(_6660_), .B(decoded_rs2_1_bF_buf16_), .C(decoded_rs2_0_bF_buf64_), .Y(_6661_) );
AOI21X1 AOI21X1_176 ( .A(decoded_rs2_1_bF_buf15_), .B(cpuregs_15_[17]), .C(_6661_), .Y(_6662_) );
AND2X2 AND2X2_34 ( .A(decoded_rs2_1_bF_buf14_), .B(cpuregs_14_[17]), .Y(_6663_) );
INVX1 INVX1_474 ( .A(cpuregs_12_[17]), .Y(_6664_) );
OAI21X1 OAI21X1_884 ( .A(_6664_), .B(decoded_rs2_1_bF_buf13_), .C(_5362__bF_buf13), .Y(_6665_) );
OAI21X1 OAI21X1_885 ( .A(_6665_), .B(_6663_), .C(decoded_rs2_2_bF_buf4_), .Y(_6666_) );
OAI22X1 OAI22X1_51 ( .A(_6659_), .B(_6655_), .C(_6662_), .D(_6666_), .Y(_6667_) );
MUX2X1 MUX2X1_102 ( .A(_6652_), .B(_6667_), .S(decoded_rs2_4_bF_buf6_), .Y(_6668_) );
NOR2X1 NOR2X1_382 ( .A(_5348__bF_buf0), .B(_6668_), .Y(_6669_) );
OAI21X1 OAI21X1_886 ( .A(_6637_), .B(_6669_), .C(_6422_), .Y(_6670_) );
AOI21X1 AOI21X1_177 ( .A(decoded_imm_17_), .B(_5849__bF_buf2), .C(_4540__bF_buf5), .Y(_6671_) );
AOI22X1 AOI22X1_26 ( .A(_5058_), .B(_4540__bF_buf4), .C(_6670_), .D(_6671_), .Y(_82__17_) );
INVX1 INVX1_475 ( .A(cpuregs_20_[18]), .Y(_6672_) );
OAI21X1 OAI21X1_887 ( .A(_5358__bF_buf4), .B(_6672_), .C(_5362__bF_buf12), .Y(_6673_) );
AOI21X1 AOI21X1_178 ( .A(_5358__bF_buf3), .B(cpuregs_16_[18]), .C(_6673_), .Y(_6674_) );
INVX1 INVX1_476 ( .A(cpuregs_21_[18]), .Y(_6675_) );
OAI21X1 OAI21X1_888 ( .A(_5358__bF_buf2), .B(_6675_), .C(decoded_rs2_0_bF_buf63_), .Y(_6676_) );
AOI21X1 AOI21X1_179 ( .A(_5358__bF_buf1), .B(cpuregs_17_[18]), .C(_6676_), .Y(_6677_) );
OAI21X1 OAI21X1_889 ( .A(_6674_), .B(_6677_), .C(_5349__bF_buf2), .Y(_6678_) );
INVX1 INVX1_477 ( .A(cpuregs_22_[18]), .Y(_6679_) );
OAI21X1 OAI21X1_890 ( .A(_5358__bF_buf0), .B(_6679_), .C(_5362__bF_buf11), .Y(_6680_) );
AOI21X1 AOI21X1_180 ( .A(_5358__bF_buf12), .B(cpuregs_18_[18]), .C(_6680_), .Y(_6681_) );
INVX1 INVX1_478 ( .A(cpuregs_23_[18]), .Y(_6682_) );
OAI21X1 OAI21X1_891 ( .A(_5358__bF_buf11), .B(_6682_), .C(decoded_rs2_0_bF_buf62_), .Y(_6683_) );
AOI21X1 AOI21X1_181 ( .A(_5358__bF_buf10), .B(cpuregs_19_[18]), .C(_6683_), .Y(_6684_) );
OAI21X1 OAI21X1_892 ( .A(_6681_), .B(_6684_), .C(decoded_rs2_1_bF_buf12_), .Y(_6685_) );
NAND3X1 NAND3X1_26 ( .A(decoded_rs2_4_bF_buf5_), .B(_6678_), .C(_6685_), .Y(_6686_) );
INVX1 INVX1_479 ( .A(cpuregs_6_[18]), .Y(_6687_) );
AOI21X1 AOI21X1_182 ( .A(decoded_rs2_1_bF_buf11_), .B(_6687_), .C(decoded_rs2_0_bF_buf61_), .Y(_6688_) );
OAI21X1 OAI21X1_893 ( .A(decoded_rs2_1_bF_buf10_), .B(cpuregs_4_[18]), .C(_6688_), .Y(_6689_) );
NOR2X1 NOR2X1_383 ( .A(cpuregs_5_[18]), .B(decoded_rs2_1_bF_buf9_), .Y(_6690_) );
OAI21X1 OAI21X1_894 ( .A(_5349__bF_buf1), .B(cpuregs_7_[18]), .C(decoded_rs2_0_bF_buf60_), .Y(_6691_) );
OAI21X1 OAI21X1_895 ( .A(_6690_), .B(_6691_), .C(_6689_), .Y(_6692_) );
INVX1 INVX1_480 ( .A(cpuregs_2_[18]), .Y(_6693_) );
AOI21X1 AOI21X1_183 ( .A(decoded_rs2_1_bF_buf8_), .B(_6693_), .C(decoded_rs2_0_bF_buf59_), .Y(_6694_) );
OAI21X1 OAI21X1_896 ( .A(decoded_rs2_1_bF_buf7_), .B(cpuregs_0_[18]), .C(_6694_), .Y(_6695_) );
NOR2X1 NOR2X1_384 ( .A(decoded_rs2_1_bF_buf6_), .B(cpuregs_1_[18]), .Y(_6696_) );
OAI21X1 OAI21X1_897 ( .A(_5349__bF_buf0), .B(cpuregs_3_[18]), .C(decoded_rs2_0_bF_buf58_), .Y(_6697_) );
OAI21X1 OAI21X1_898 ( .A(_6696_), .B(_6697_), .C(_6695_), .Y(_6698_) );
MUX2X1 MUX2X1_103 ( .A(_6698_), .B(_6692_), .S(_5358__bF_buf9), .Y(_6699_) );
OAI21X1 OAI21X1_899 ( .A(decoded_rs2_4_bF_buf4_), .B(_6699_), .C(_6686_), .Y(_6700_) );
AND2X2 AND2X2_35 ( .A(_6700_), .B(_5348__bF_buf5), .Y(_6701_) );
INVX1 INVX1_481 ( .A(cpuregs_28_[18]), .Y(_6702_) );
NAND2X1 NAND2X1_388 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_29_[18]), .Y(_6703_) );
OAI21X1 OAI21X1_900 ( .A(_6702_), .B(decoded_rs2_0_bF_buf56_), .C(_6703_), .Y(_6704_) );
INVX1 INVX1_482 ( .A(cpuregs_31_[18]), .Y(_6705_) );
OAI21X1 OAI21X1_901 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_30_[18]), .C(decoded_rs2_1_bF_buf5_), .Y(_6706_) );
AOI21X1 AOI21X1_184 ( .A(decoded_rs2_0_bF_buf54_), .B(_6705_), .C(_6706_), .Y(_6707_) );
AOI21X1 AOI21X1_185 ( .A(_5349__bF_buf11), .B(_6704_), .C(_6707_), .Y(_6708_) );
NOR2X1 NOR2X1_385 ( .A(_5358__bF_buf8), .B(_6708_), .Y(_6709_) );
INVX1 INVX1_483 ( .A(cpuregs_24_[18]), .Y(_6710_) );
NAND2X1 NAND2X1_389 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_25_[18]), .Y(_6711_) );
OAI21X1 OAI21X1_902 ( .A(_6710_), .B(decoded_rs2_0_bF_buf52_), .C(_6711_), .Y(_6712_) );
INVX1 INVX1_484 ( .A(cpuregs_27_[18]), .Y(_6713_) );
OAI21X1 OAI21X1_903 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_26_[18]), .C(decoded_rs2_1_bF_buf4_), .Y(_6714_) );
AOI21X1 AOI21X1_186 ( .A(decoded_rs2_0_bF_buf50_), .B(_6713_), .C(_6714_), .Y(_6715_) );
AOI21X1 AOI21X1_187 ( .A(_5349__bF_buf10), .B(_6712_), .C(_6715_), .Y(_6716_) );
NOR2X1 NOR2X1_386 ( .A(decoded_rs2_2_bF_buf3_), .B(_6716_), .Y(_6717_) );
OAI21X1 OAI21X1_904 ( .A(_6709_), .B(_6717_), .C(decoded_rs2_4_bF_buf3_), .Y(_6718_) );
NOR2X1 NOR2X1_387 ( .A(cpuregs_8_[18]), .B(decoded_rs2_0_bF_buf49_), .Y(_6719_) );
OAI21X1 OAI21X1_905 ( .A(_5362__bF_buf10), .B(cpuregs_9_[18]), .C(_5349__bF_buf9), .Y(_6720_) );
NOR2X1 NOR2X1_388 ( .A(cpuregs_11_[18]), .B(_5362__bF_buf9), .Y(_6721_) );
OAI21X1 OAI21X1_906 ( .A(decoded_rs2_0_bF_buf48_), .B(cpuregs_10_[18]), .C(decoded_rs2_1_bF_buf3_), .Y(_6722_) );
OAI22X1 OAI22X1_52 ( .A(_6721_), .B(_6722_), .C(_6720_), .D(_6719_), .Y(_6723_) );
INVX1 INVX1_485 ( .A(cpuregs_13_[18]), .Y(_6724_) );
AOI21X1 AOI21X1_188 ( .A(decoded_rs2_0_bF_buf47_), .B(_6724_), .C(decoded_rs2_1_bF_buf2_), .Y(_6725_) );
OAI21X1 OAI21X1_907 ( .A(decoded_rs2_0_bF_buf46_), .B(cpuregs_12_[18]), .C(_6725_), .Y(_6726_) );
NOR2X1 NOR2X1_389 ( .A(cpuregs_15_[18]), .B(_5362__bF_buf8), .Y(_6727_) );
OAI21X1 OAI21X1_908 ( .A(decoded_rs2_0_bF_buf45_), .B(cpuregs_14_[18]), .C(decoded_rs2_1_bF_buf1_), .Y(_6728_) );
OAI21X1 OAI21X1_909 ( .A(_6727_), .B(_6728_), .C(_6726_), .Y(_6729_) );
MUX2X1 MUX2X1_104 ( .A(_6729_), .B(_6723_), .S(decoded_rs2_2_bF_buf2_), .Y(_6730_) );
OAI21X1 OAI21X1_910 ( .A(decoded_rs2_4_bF_buf2_), .B(_6730_), .C(_6718_), .Y(_6731_) );
AND2X2 AND2X2_36 ( .A(_6731_), .B(decoded_rs2_3_bF_buf2_), .Y(_6732_) );
OAI21X1 OAI21X1_911 ( .A(_6732_), .B(_6701_), .C(_6422_), .Y(_6733_) );
AOI21X1 AOI21X1_189 ( .A(decoded_imm_18_), .B(_5849__bF_buf1), .C(_4540__bF_buf3), .Y(_6734_) );
AOI22X1 AOI22X1_27 ( .A(_5046_), .B(_4540__bF_buf2), .C(_6733_), .D(_6734_), .Y(_82__18_) );
INVX1 INVX1_486 ( .A(cpuregs_28_[19]), .Y(_6735_) );
OAI21X1 OAI21X1_912 ( .A(_5358__bF_buf7), .B(_6735_), .C(_5362__bF_buf7), .Y(_6736_) );
AOI21X1 AOI21X1_190 ( .A(_5358__bF_buf6), .B(cpuregs_24_[19]), .C(_6736_), .Y(_6737_) );
INVX1 INVX1_487 ( .A(cpuregs_29_[19]), .Y(_6738_) );
OAI21X1 OAI21X1_913 ( .A(_5358__bF_buf5), .B(_6738_), .C(decoded_rs2_0_bF_buf44_), .Y(_6739_) );
AOI21X1 AOI21X1_191 ( .A(_5358__bF_buf4), .B(cpuregs_25_[19]), .C(_6739_), .Y(_6740_) );
OAI21X1 OAI21X1_914 ( .A(_6737_), .B(_6740_), .C(_5349__bF_buf8), .Y(_6741_) );
INVX1 INVX1_488 ( .A(cpuregs_30_[19]), .Y(_6742_) );
OAI21X1 OAI21X1_915 ( .A(_5358__bF_buf3), .B(_6742_), .C(_5362__bF_buf6), .Y(_6743_) );
AOI21X1 AOI21X1_192 ( .A(_5358__bF_buf2), .B(cpuregs_26_[19]), .C(_6743_), .Y(_6744_) );
INVX1 INVX1_489 ( .A(cpuregs_31_[19]), .Y(_6745_) );
OAI21X1 OAI21X1_916 ( .A(_5358__bF_buf1), .B(_6745_), .C(decoded_rs2_0_bF_buf43_), .Y(_6746_) );
AOI21X1 AOI21X1_193 ( .A(_5358__bF_buf0), .B(cpuregs_27_[19]), .C(_6746_), .Y(_6747_) );
OAI21X1 OAI21X1_917 ( .A(_6744_), .B(_6747_), .C(decoded_rs2_1_bF_buf0_), .Y(_6748_) );
NAND3X1 NAND3X1_27 ( .A(decoded_rs2_4_bF_buf1_), .B(_6741_), .C(_6748_), .Y(_6749_) );
NOR2X1 NOR2X1_390 ( .A(cpuregs_8_[19]), .B(decoded_rs2_0_bF_buf42_), .Y(_6750_) );
OAI21X1 OAI21X1_918 ( .A(_5362__bF_buf5), .B(cpuregs_9_[19]), .C(_5349__bF_buf7), .Y(_6751_) );
NOR2X1 NOR2X1_391 ( .A(cpuregs_11_[19]), .B(_5362__bF_buf4), .Y(_6752_) );
OAI21X1 OAI21X1_919 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_10_[19]), .C(decoded_rs2_1_bF_buf45_), .Y(_6753_) );
OAI22X1 OAI22X1_53 ( .A(_6752_), .B(_6753_), .C(_6751_), .D(_6750_), .Y(_6754_) );
INVX1 INVX1_490 ( .A(cpuregs_13_[19]), .Y(_6755_) );
AOI21X1 AOI21X1_194 ( .A(decoded_rs2_0_bF_buf40_), .B(_6755_), .C(decoded_rs2_1_bF_buf44_), .Y(_6756_) );
OAI21X1 OAI21X1_920 ( .A(decoded_rs2_0_bF_buf39_), .B(cpuregs_12_[19]), .C(_6756_), .Y(_6757_) );
NOR2X1 NOR2X1_392 ( .A(cpuregs_15_[19]), .B(_5362__bF_buf3), .Y(_6758_) );
OAI21X1 OAI21X1_921 ( .A(decoded_rs2_0_bF_buf38_), .B(cpuregs_14_[19]), .C(decoded_rs2_1_bF_buf43_), .Y(_6759_) );
OAI21X1 OAI21X1_922 ( .A(_6758_), .B(_6759_), .C(_6757_), .Y(_6760_) );
MUX2X1 MUX2X1_105 ( .A(_6760_), .B(_6754_), .S(decoded_rs2_2_bF_buf1_), .Y(_6761_) );
OAI21X1 OAI21X1_923 ( .A(decoded_rs2_4_bF_buf0_), .B(_6761_), .C(_6749_), .Y(_6762_) );
AND2X2 AND2X2_37 ( .A(_6762_), .B(decoded_rs2_3_bF_buf1_), .Y(_6763_) );
INVX1 INVX1_491 ( .A(cpuregs_17_[19]), .Y(_6764_) );
AOI21X1 AOI21X1_195 ( .A(decoded_rs2_0_bF_buf37_), .B(_6764_), .C(decoded_rs2_1_bF_buf42_), .Y(_6765_) );
OAI21X1 OAI21X1_924 ( .A(decoded_rs2_0_bF_buf36_), .B(cpuregs_16_[19]), .C(_6765_), .Y(_6766_) );
NOR2X1 NOR2X1_393 ( .A(cpuregs_19_[19]), .B(_5362__bF_buf2), .Y(_6767_) );
OAI21X1 OAI21X1_925 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_18_[19]), .C(decoded_rs2_1_bF_buf41_), .Y(_6768_) );
OAI21X1 OAI21X1_926 ( .A(_6767_), .B(_6768_), .C(_6766_), .Y(_6769_) );
INVX1 INVX1_492 ( .A(cpuregs_20_[19]), .Y(_6770_) );
NAND2X1 NAND2X1_390 ( .A(decoded_rs2_0_bF_buf34_), .B(cpuregs_21_[19]), .Y(_6771_) );
OAI21X1 OAI21X1_927 ( .A(_6770_), .B(decoded_rs2_0_bF_buf33_), .C(_6771_), .Y(_6772_) );
INVX1 INVX1_493 ( .A(cpuregs_22_[19]), .Y(_6773_) );
NAND2X1 NAND2X1_391 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_23_[19]), .Y(_6774_) );
OAI21X1 OAI21X1_928 ( .A(_6773_), .B(decoded_rs2_0_bF_buf31_), .C(_6774_), .Y(_6775_) );
MUX2X1 MUX2X1_106 ( .A(_6775_), .B(_6772_), .S(decoded_rs2_1_bF_buf40_), .Y(_6776_) );
NOR2X1 NOR2X1_394 ( .A(_5358__bF_buf12), .B(_6776_), .Y(_6777_) );
AOI21X1 AOI21X1_196 ( .A(_5358__bF_buf11), .B(_6769_), .C(_6777_), .Y(_6778_) );
NOR2X1 NOR2X1_395 ( .A(decoded_rs2_0_bF_buf30_), .B(cpuregs_4_[19]), .Y(_6779_) );
OAI21X1 OAI21X1_929 ( .A(_5362__bF_buf1), .B(cpuregs_5_[19]), .C(_5349__bF_buf6), .Y(_6780_) );
NOR2X1 NOR2X1_396 ( .A(cpuregs_7_[19]), .B(_5362__bF_buf0), .Y(_6781_) );
OAI21X1 OAI21X1_930 ( .A(cpuregs_6_[19]), .B(decoded_rs2_0_bF_buf29_), .C(decoded_rs2_1_bF_buf39_), .Y(_6782_) );
OAI22X1 OAI22X1_54 ( .A(_6781_), .B(_6782_), .C(_6780_), .D(_6779_), .Y(_6783_) );
NOR2X1 NOR2X1_397 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_0_[19]), .Y(_6784_) );
OAI21X1 OAI21X1_931 ( .A(_5362__bF_buf14), .B(cpuregs_1_[19]), .C(_5349__bF_buf5), .Y(_6785_) );
NOR2X1 NOR2X1_398 ( .A(cpuregs_3_[19]), .B(_5362__bF_buf13), .Y(_6786_) );
OAI21X1 OAI21X1_932 ( .A(decoded_rs2_0_bF_buf27_), .B(cpuregs_2_[19]), .C(decoded_rs2_1_bF_buf38_), .Y(_6787_) );
OAI22X1 OAI22X1_55 ( .A(_6786_), .B(_6787_), .C(_6785_), .D(_6784_), .Y(_6788_) );
MUX2X1 MUX2X1_107 ( .A(_6788_), .B(_6783_), .S(_5358__bF_buf10), .Y(_6789_) );
MUX2X1 MUX2X1_108 ( .A(_6778_), .B(_6789_), .S(decoded_rs2_4_bF_buf7_), .Y(_6790_) );
AND2X2 AND2X2_38 ( .A(_6790_), .B(_5348__bF_buf4), .Y(_6791_) );
OAI21X1 OAI21X1_933 ( .A(_6791_), .B(_6763_), .C(_6422_), .Y(_6792_) );
AOI21X1 AOI21X1_197 ( .A(decoded_imm_19_), .B(_5849__bF_buf0), .C(_4540__bF_buf1), .Y(_6793_) );
AOI22X1 AOI22X1_28 ( .A(_5041_), .B(_4540__bF_buf0), .C(_6792_), .D(_6793_), .Y(_82__19_) );
NOR2X1 NOR2X1_399 ( .A(_10735__20_), .B(_4539__bF_buf0), .Y(_6794_) );
INVX1 INVX1_494 ( .A(cpuregs_24_[20]), .Y(_6795_) );
NAND2X1 NAND2X1_392 ( .A(decoded_rs2_1_bF_buf37_), .B(cpuregs_26_[20]), .Y(_6796_) );
OAI21X1 OAI21X1_934 ( .A(_6795_), .B(decoded_rs2_1_bF_buf36_), .C(_6796_), .Y(_6797_) );
MUX2X1 MUX2X1_109 ( .A(cpuregs_27_[20]), .B(cpuregs_25_[20]), .S(decoded_rs2_1_bF_buf35_), .Y(_6798_) );
OAI21X1 OAI21X1_935 ( .A(_6798_), .B(_5362__bF_buf12), .C(_5358__bF_buf9), .Y(_6799_) );
AOI21X1 AOI21X1_198 ( .A(_5362__bF_buf11), .B(_6797_), .C(_6799_), .Y(_6800_) );
NOR2X1 NOR2X1_400 ( .A(decoded_rs2_0_bF_buf26_), .B(cpuregs_28_[20]), .Y(_6801_) );
OAI21X1 OAI21X1_936 ( .A(_5362__bF_buf10), .B(cpuregs_29_[20]), .C(_5349__bF_buf4), .Y(_6802_) );
NOR2X1 NOR2X1_401 ( .A(cpuregs_31_[20]), .B(_5362__bF_buf9), .Y(_6803_) );
OAI21X1 OAI21X1_937 ( .A(decoded_rs2_0_bF_buf25_), .B(cpuregs_30_[20]), .C(decoded_rs2_1_bF_buf34_), .Y(_6804_) );
OAI22X1 OAI22X1_56 ( .A(_6803_), .B(_6804_), .C(_6802_), .D(_6801_), .Y(_6805_) );
OAI21X1 OAI21X1_938 ( .A(_6805_), .B(_5358__bF_buf8), .C(decoded_rs2_3_bF_buf0_), .Y(_6806_) );
INVX1 INVX1_495 ( .A(cpuregs_17_[20]), .Y(_6807_) );
AOI21X1 AOI21X1_199 ( .A(decoded_rs2_0_bF_buf24_), .B(_6807_), .C(decoded_rs2_1_bF_buf33_), .Y(_6808_) );
OAI21X1 OAI21X1_939 ( .A(decoded_rs2_0_bF_buf23_), .B(cpuregs_16_[20]), .C(_6808_), .Y(_6809_) );
INVX1 INVX1_496 ( .A(cpuregs_18_[20]), .Y(_6810_) );
AOI21X1 AOI21X1_200 ( .A(_5362__bF_buf8), .B(_6810_), .C(_5349__bF_buf3), .Y(_6811_) );
OAI21X1 OAI21X1_940 ( .A(_5362__bF_buf7), .B(cpuregs_19_[20]), .C(_6811_), .Y(_6812_) );
NAND3X1 NAND3X1_28 ( .A(_5358__bF_buf7), .B(_6809_), .C(_6812_), .Y(_6813_) );
INVX1 INVX1_497 ( .A(cpuregs_21_[20]), .Y(_6814_) );
AOI21X1 AOI21X1_201 ( .A(decoded_rs2_0_bF_buf22_), .B(_6814_), .C(decoded_rs2_1_bF_buf32_), .Y(_6815_) );
OAI21X1 OAI21X1_941 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_20_[20]), .C(_6815_), .Y(_6816_) );
NOR2X1 NOR2X1_402 ( .A(cpuregs_23_[20]), .B(_5362__bF_buf6), .Y(_6817_) );
OAI21X1 OAI21X1_942 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_22_[20]), .C(decoded_rs2_1_bF_buf31_), .Y(_6818_) );
OAI21X1 OAI21X1_943 ( .A(_6817_), .B(_6818_), .C(_6816_), .Y(_6819_) );
OAI21X1 OAI21X1_944 ( .A(_6819_), .B(_5358__bF_buf6), .C(_6813_), .Y(_6820_) );
OAI22X1 OAI22X1_57 ( .A(_6800_), .B(_6806_), .C(_6820_), .D(decoded_rs2_3_bF_buf6_), .Y(_6821_) );
NAND2X1 NAND2X1_393 ( .A(decoded_rs2_4_bF_buf6_), .B(_6821_), .Y(_6822_) );
INVX1 INVX1_498 ( .A(cpuregs_8_[20]), .Y(_6823_) );
OAI21X1 OAI21X1_945 ( .A(_5362__bF_buf5), .B(cpuregs_9_[20]), .C(_5349__bF_buf2), .Y(_6824_) );
AOI21X1 AOI21X1_202 ( .A(_6823_), .B(_5362__bF_buf4), .C(_6824_), .Y(_6825_) );
INVX1 INVX1_499 ( .A(cpuregs_11_[20]), .Y(_6826_) );
OAI21X1 OAI21X1_946 ( .A(decoded_rs2_0_bF_buf19_), .B(cpuregs_10_[20]), .C(decoded_rs2_1_bF_buf30_), .Y(_6827_) );
AOI21X1 AOI21X1_203 ( .A(decoded_rs2_0_bF_buf18_), .B(_6826_), .C(_6827_), .Y(_6828_) );
OAI21X1 OAI21X1_947 ( .A(_6825_), .B(_6828_), .C(_5358__bF_buf5), .Y(_6829_) );
INVX1 INVX1_500 ( .A(cpuregs_12_[20]), .Y(_6830_) );
OAI21X1 OAI21X1_948 ( .A(_5362__bF_buf3), .B(cpuregs_13_[20]), .C(_5349__bF_buf1), .Y(_6831_) );
AOI21X1 AOI21X1_204 ( .A(_5362__bF_buf2), .B(_6830_), .C(_6831_), .Y(_6832_) );
INVX1 INVX1_501 ( .A(cpuregs_15_[20]), .Y(_6833_) );
OAI21X1 OAI21X1_949 ( .A(decoded_rs2_0_bF_buf17_), .B(cpuregs_14_[20]), .C(decoded_rs2_1_bF_buf29_), .Y(_6834_) );
AOI21X1 AOI21X1_205 ( .A(decoded_rs2_0_bF_buf16_), .B(_6833_), .C(_6834_), .Y(_6835_) );
OAI21X1 OAI21X1_950 ( .A(_6832_), .B(_6835_), .C(decoded_rs2_2_bF_buf0_), .Y(_6836_) );
AOI21X1 AOI21X1_206 ( .A(_6829_), .B(_6836_), .C(_5348__bF_buf3), .Y(_6837_) );
NOR2X1 NOR2X1_403 ( .A(decoded_rs2_0_bF_buf15_), .B(cpuregs_0_[20]), .Y(_6838_) );
OAI21X1 OAI21X1_951 ( .A(_5362__bF_buf1), .B(cpuregs_1_[20]), .C(_5349__bF_buf0), .Y(_6839_) );
NOR2X1 NOR2X1_404 ( .A(cpuregs_3_[20]), .B(_5362__bF_buf0), .Y(_6840_) );
OAI21X1 OAI21X1_952 ( .A(decoded_rs2_0_bF_buf14_), .B(cpuregs_2_[20]), .C(decoded_rs2_1_bF_buf28_), .Y(_6841_) );
OAI22X1 OAI22X1_58 ( .A(_6840_), .B(_6841_), .C(_6839_), .D(_6838_), .Y(_6842_) );
NAND2X1 NAND2X1_394 ( .A(_5358__bF_buf4), .B(_6842_), .Y(_6843_) );
INVX1 INVX1_502 ( .A(cpuregs_4_[20]), .Y(_6844_) );
NAND2X1 NAND2X1_395 ( .A(cpuregs_5_[20]), .B(decoded_rs2_0_bF_buf13_), .Y(_6845_) );
OAI21X1 OAI21X1_953 ( .A(_6844_), .B(decoded_rs2_0_bF_buf12_), .C(_6845_), .Y(_6846_) );
INVX1 INVX1_503 ( .A(cpuregs_6_[20]), .Y(_6847_) );
NAND2X1 NAND2X1_396 ( .A(cpuregs_7_[20]), .B(decoded_rs2_0_bF_buf11_), .Y(_6848_) );
OAI21X1 OAI21X1_954 ( .A(_6847_), .B(decoded_rs2_0_bF_buf10_), .C(_6848_), .Y(_6849_) );
MUX2X1 MUX2X1_110 ( .A(_6849_), .B(_6846_), .S(decoded_rs2_1_bF_buf27_), .Y(_6850_) );
OAI21X1 OAI21X1_955 ( .A(_5358__bF_buf3), .B(_6850_), .C(_6843_), .Y(_6851_) );
AOI21X1 AOI21X1_207 ( .A(_5348__bF_buf2), .B(_6851_), .C(_6837_), .Y(_6852_) );
OAI21X1 OAI21X1_956 ( .A(decoded_rs2_4_bF_buf5_), .B(_6852_), .C(_6822_), .Y(_6853_) );
NAND2X1 NAND2X1_397 ( .A(_6422_), .B(_6853_), .Y(_6854_) );
AOI21X1 AOI21X1_208 ( .A(decoded_imm_20_), .B(_5849__bF_buf4), .C(_4540__bF_buf6), .Y(_6855_) );
AOI21X1 AOI21X1_209 ( .A(_6855_), .B(_6854_), .C(_6794_), .Y(_82__20_) );
NOR2X1 NOR2X1_405 ( .A(_10735__21_), .B(_4539__bF_buf3), .Y(_6856_) );
NOR2X1 NOR2X1_406 ( .A(decoded_rs2_0_bF_buf9_), .B(cpuregs_0_[21]), .Y(_6857_) );
OAI21X1 OAI21X1_957 ( .A(_5362__bF_buf14), .B(cpuregs_1_[21]), .C(_5349__bF_buf11), .Y(_6858_) );
NOR2X1 NOR2X1_407 ( .A(cpuregs_3_[21]), .B(_5362__bF_buf13), .Y(_6859_) );
OAI21X1 OAI21X1_958 ( .A(decoded_rs2_0_bF_buf8_), .B(cpuregs_2_[21]), .C(decoded_rs2_1_bF_buf26_), .Y(_6860_) );
OAI22X1 OAI22X1_59 ( .A(_6859_), .B(_6860_), .C(_6858_), .D(_6857_), .Y(_6861_) );
NOR2X1 NOR2X1_408 ( .A(decoded_rs2_2_bF_buf8_), .B(_6861_), .Y(_6862_) );
NOR2X1 NOR2X1_409 ( .A(decoded_rs2_0_bF_buf7_), .B(cpuregs_4_[21]), .Y(_6863_) );
OAI21X1 OAI21X1_959 ( .A(_5362__bF_buf12), .B(cpuregs_5_[21]), .C(_5349__bF_buf10), .Y(_6864_) );
NOR2X1 NOR2X1_410 ( .A(cpuregs_7_[21]), .B(_5362__bF_buf11), .Y(_6865_) );
OAI21X1 OAI21X1_960 ( .A(cpuregs_6_[21]), .B(decoded_rs2_0_bF_buf6_), .C(decoded_rs2_1_bF_buf25_), .Y(_6866_) );
OAI22X1 OAI22X1_60 ( .A(_6865_), .B(_6866_), .C(_6864_), .D(_6863_), .Y(_6867_) );
OAI21X1 OAI21X1_961 ( .A(_6867_), .B(_5358__bF_buf2), .C(_5348__bF_buf1), .Y(_6868_) );
NOR2X1 NOR2X1_411 ( .A(decoded_rs2_0_bF_buf5_), .B(cpuregs_12_[21]), .Y(_6869_) );
OAI21X1 OAI21X1_962 ( .A(_5362__bF_buf10), .B(cpuregs_13_[21]), .C(_5349__bF_buf9), .Y(_6870_) );
NOR2X1 NOR2X1_412 ( .A(cpuregs_15_[21]), .B(_5362__bF_buf9), .Y(_6871_) );
OAI21X1 OAI21X1_963 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_14_[21]), .C(decoded_rs2_1_bF_buf24_), .Y(_6872_) );
OAI22X1 OAI22X1_61 ( .A(_6871_), .B(_6872_), .C(_6870_), .D(_6869_), .Y(_6873_) );
NOR2X1 NOR2X1_413 ( .A(_5358__bF_buf1), .B(_6873_), .Y(_6874_) );
NOR2X1 NOR2X1_414 ( .A(cpuregs_8_[21]), .B(decoded_rs2_0_bF_buf3_), .Y(_6875_) );
OAI21X1 OAI21X1_964 ( .A(_5362__bF_buf8), .B(cpuregs_9_[21]), .C(_5349__bF_buf8), .Y(_6876_) );
NOR2X1 NOR2X1_415 ( .A(cpuregs_11_[21]), .B(_5362__bF_buf7), .Y(_6877_) );
OAI21X1 OAI21X1_965 ( .A(decoded_rs2_0_bF_buf2_), .B(cpuregs_10_[21]), .C(decoded_rs2_1_bF_buf23_), .Y(_6878_) );
OAI22X1 OAI22X1_62 ( .A(_6877_), .B(_6878_), .C(_6876_), .D(_6875_), .Y(_6879_) );
OAI21X1 OAI21X1_966 ( .A(_6879_), .B(decoded_rs2_2_bF_buf7_), .C(decoded_rs2_3_bF_buf5_), .Y(_6880_) );
OAI22X1 OAI22X1_63 ( .A(_6868_), .B(_6862_), .C(_6874_), .D(_6880_), .Y(_6881_) );
INVX1 INVX1_504 ( .A(cpuregs_26_[21]), .Y(_6882_) );
OAI21X1 OAI21X1_967 ( .A(_6882_), .B(decoded_rs2_0_bF_buf1_), .C(decoded_rs2_1_bF_buf22_), .Y(_6883_) );
AOI21X1 AOI21X1_210 ( .A(decoded_rs2_0_bF_buf0_), .B(cpuregs_27_[21]), .C(_6883_), .Y(_6884_) );
AND2X2 AND2X2_39 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_25_[21]), .Y(_6885_) );
INVX1 INVX1_505 ( .A(cpuregs_24_[21]), .Y(_6886_) );
OAI21X1 OAI21X1_968 ( .A(_6886_), .B(decoded_rs2_0_bF_buf77_), .C(_5349__bF_buf7), .Y(_6887_) );
OAI21X1 OAI21X1_969 ( .A(_6887_), .B(_6885_), .C(_5358__bF_buf0), .Y(_6888_) );
INVX1 INVX1_506 ( .A(cpuregs_28_[21]), .Y(_6889_) );
NAND2X1 NAND2X1_398 ( .A(decoded_rs2_0_bF_buf76_), .B(cpuregs_29_[21]), .Y(_6890_) );
OAI21X1 OAI21X1_970 ( .A(_6889_), .B(decoded_rs2_0_bF_buf75_), .C(_6890_), .Y(_6891_) );
INVX1 INVX1_507 ( .A(cpuregs_30_[21]), .Y(_6892_) );
NAND2X1 NAND2X1_399 ( .A(decoded_rs2_0_bF_buf74_), .B(cpuregs_31_[21]), .Y(_6893_) );
OAI21X1 OAI21X1_971 ( .A(_6892_), .B(decoded_rs2_0_bF_buf73_), .C(_6893_), .Y(_6894_) );
MUX2X1 MUX2X1_111 ( .A(_6894_), .B(_6891_), .S(decoded_rs2_1_bF_buf21_), .Y(_6895_) );
OAI22X1 OAI22X1_64 ( .A(_6888_), .B(_6884_), .C(_6895_), .D(_5358__bF_buf12), .Y(_6896_) );
INVX1 INVX1_508 ( .A(cpuregs_16_[21]), .Y(_6897_) );
NAND2X1 NAND2X1_400 ( .A(decoded_rs2_0_bF_buf72_), .B(cpuregs_17_[21]), .Y(_6898_) );
OAI21X1 OAI21X1_972 ( .A(_6897_), .B(decoded_rs2_0_bF_buf71_), .C(_6898_), .Y(_6899_) );
INVX1 INVX1_509 ( .A(cpuregs_19_[21]), .Y(_6900_) );
OAI21X1 OAI21X1_973 ( .A(decoded_rs2_0_bF_buf70_), .B(cpuregs_18_[21]), .C(decoded_rs2_1_bF_buf20_), .Y(_6901_) );
AOI21X1 AOI21X1_211 ( .A(decoded_rs2_0_bF_buf69_), .B(_6900_), .C(_6901_), .Y(_6902_) );
AOI21X1 AOI21X1_212 ( .A(_5349__bF_buf6), .B(_6899_), .C(_6902_), .Y(_6903_) );
NAND2X1 NAND2X1_401 ( .A(_5358__bF_buf11), .B(_6903_), .Y(_6904_) );
INVX1 INVX1_510 ( .A(cpuregs_21_[21]), .Y(_6905_) );
NAND2X1 NAND2X1_402 ( .A(cpuregs_20_[21]), .B(_5362__bF_buf6), .Y(_6906_) );
OAI21X1 OAI21X1_974 ( .A(_5362__bF_buf5), .B(_6905_), .C(_6906_), .Y(_6907_) );
INVX1 INVX1_511 ( .A(cpuregs_22_[21]), .Y(_6908_) );
NAND2X1 NAND2X1_403 ( .A(decoded_rs2_0_bF_buf68_), .B(cpuregs_23_[21]), .Y(_6909_) );
OAI21X1 OAI21X1_975 ( .A(_6908_), .B(decoded_rs2_0_bF_buf67_), .C(_6909_), .Y(_6910_) );
MUX2X1 MUX2X1_112 ( .A(_6907_), .B(_6910_), .S(_5349__bF_buf5), .Y(_6911_) );
AOI21X1 AOI21X1_213 ( .A(decoded_rs2_2_bF_buf6_), .B(_6911_), .C(decoded_rs2_3_bF_buf4_), .Y(_6912_) );
AOI22X1 AOI22X1_29 ( .A(decoded_rs2_3_bF_buf3_), .B(_6896_), .C(_6912_), .D(_6904_), .Y(_6913_) );
AOI21X1 AOI21X1_214 ( .A(decoded_rs2_4_bF_buf4_), .B(_6913_), .C(_5890__bF_buf0), .Y(_6914_) );
OAI21X1 OAI21X1_976 ( .A(decoded_rs2_4_bF_buf3_), .B(_6881_), .C(_6914_), .Y(_6915_) );
AOI21X1 AOI21X1_215 ( .A(decoded_imm_21_), .B(_5849__bF_buf3), .C(_4540__bF_buf5), .Y(_6916_) );
AOI21X1 AOI21X1_216 ( .A(_6916_), .B(_6915_), .C(_6856_), .Y(_82__21_) );
NOR2X1 NOR2X1_416 ( .A(decoded_rs2_0_bF_buf66_), .B(cpuregs_4_[22]), .Y(_6917_) );
OAI21X1 OAI21X1_977 ( .A(_5362__bF_buf4), .B(cpuregs_5_[22]), .C(_5349__bF_buf4), .Y(_6918_) );
NOR2X1 NOR2X1_417 ( .A(cpuregs_7_[22]), .B(_5362__bF_buf3), .Y(_6919_) );
OAI21X1 OAI21X1_978 ( .A(cpuregs_6_[22]), .B(decoded_rs2_0_bF_buf65_), .C(decoded_rs2_1_bF_buf19_), .Y(_6920_) );
OAI22X1 OAI22X1_65 ( .A(_6919_), .B(_6920_), .C(_6918_), .D(_6917_), .Y(_6921_) );
INVX1 INVX1_512 ( .A(cpuregs_2_[22]), .Y(_6922_) );
AOI21X1 AOI21X1_217 ( .A(decoded_rs2_1_bF_buf18_), .B(_6922_), .C(decoded_rs2_0_bF_buf64_), .Y(_6923_) );
OAI21X1 OAI21X1_979 ( .A(decoded_rs2_1_bF_buf17_), .B(cpuregs_0_[22]), .C(_6923_), .Y(_6924_) );
NOR2X1 NOR2X1_418 ( .A(decoded_rs2_1_bF_buf16_), .B(cpuregs_1_[22]), .Y(_6925_) );
OAI21X1 OAI21X1_980 ( .A(_5349__bF_buf3), .B(cpuregs_3_[22]), .C(decoded_rs2_0_bF_buf63_), .Y(_6926_) );
OAI21X1 OAI21X1_981 ( .A(_6925_), .B(_6926_), .C(_6924_), .Y(_6927_) );
MUX2X1 MUX2X1_113 ( .A(_6927_), .B(_6921_), .S(_5358__bF_buf10), .Y(_6928_) );
NOR2X1 NOR2X1_419 ( .A(cpuregs_8_[22]), .B(decoded_rs2_0_bF_buf62_), .Y(_6929_) );
OAI21X1 OAI21X1_982 ( .A(_5362__bF_buf2), .B(cpuregs_9_[22]), .C(_5349__bF_buf2), .Y(_6930_) );
NOR2X1 NOR2X1_420 ( .A(cpuregs_11_[22]), .B(_5362__bF_buf1), .Y(_6931_) );
OAI21X1 OAI21X1_983 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_10_[22]), .C(decoded_rs2_1_bF_buf15_), .Y(_6932_) );
OAI22X1 OAI22X1_66 ( .A(_6931_), .B(_6932_), .C(_6930_), .D(_6929_), .Y(_6933_) );
INVX1 INVX1_513 ( .A(cpuregs_13_[22]), .Y(_6934_) );
AOI21X1 AOI21X1_218 ( .A(decoded_rs2_0_bF_buf60_), .B(_6934_), .C(decoded_rs2_1_bF_buf14_), .Y(_6935_) );
OAI21X1 OAI21X1_984 ( .A(decoded_rs2_0_bF_buf59_), .B(cpuregs_12_[22]), .C(_6935_), .Y(_6936_) );
NOR2X1 NOR2X1_421 ( .A(cpuregs_15_[22]), .B(_5362__bF_buf0), .Y(_6937_) );
OAI21X1 OAI21X1_985 ( .A(decoded_rs2_0_bF_buf58_), .B(cpuregs_14_[22]), .C(decoded_rs2_1_bF_buf13_), .Y(_6938_) );
OAI21X1 OAI21X1_986 ( .A(_6937_), .B(_6938_), .C(_6936_), .Y(_6939_) );
MUX2X1 MUX2X1_114 ( .A(_6939_), .B(_6933_), .S(decoded_rs2_2_bF_buf5_), .Y(_6940_) );
MUX2X1 MUX2X1_115 ( .A(_6940_), .B(_6928_), .S(decoded_rs2_3_bF_buf2_), .Y(_6941_) );
INVX1 INVX1_514 ( .A(cpuregs_28_[22]), .Y(_6942_) );
NAND2X1 NAND2X1_404 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_29_[22]), .Y(_6943_) );
OAI21X1 OAI21X1_987 ( .A(_6942_), .B(decoded_rs2_0_bF_buf56_), .C(_6943_), .Y(_6944_) );
INVX1 INVX1_515 ( .A(cpuregs_31_[22]), .Y(_6945_) );
OAI21X1 OAI21X1_988 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_30_[22]), .C(decoded_rs2_1_bF_buf12_), .Y(_6946_) );
AOI21X1 AOI21X1_219 ( .A(decoded_rs2_0_bF_buf54_), .B(_6945_), .C(_6946_), .Y(_6947_) );
AOI21X1 AOI21X1_220 ( .A(_5349__bF_buf1), .B(_6944_), .C(_6947_), .Y(_6948_) );
NOR2X1 NOR2X1_422 ( .A(_5358__bF_buf9), .B(_6948_), .Y(_6949_) );
INVX1 INVX1_516 ( .A(cpuregs_24_[22]), .Y(_6950_) );
NAND2X1 NAND2X1_405 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_25_[22]), .Y(_6951_) );
OAI21X1 OAI21X1_989 ( .A(_6950_), .B(decoded_rs2_0_bF_buf52_), .C(_6951_), .Y(_6952_) );
INVX1 INVX1_517 ( .A(cpuregs_27_[22]), .Y(_6953_) );
OAI21X1 OAI21X1_990 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_26_[22]), .C(decoded_rs2_1_bF_buf11_), .Y(_6954_) );
AOI21X1 AOI21X1_221 ( .A(decoded_rs2_0_bF_buf50_), .B(_6953_), .C(_6954_), .Y(_6955_) );
AOI21X1 AOI21X1_222 ( .A(_5349__bF_buf0), .B(_6952_), .C(_6955_), .Y(_6956_) );
NOR2X1 NOR2X1_423 ( .A(decoded_rs2_2_bF_buf4_), .B(_6956_), .Y(_6957_) );
OAI21X1 OAI21X1_991 ( .A(_6949_), .B(_6957_), .C(decoded_rs2_3_bF_buf1_), .Y(_6958_) );
INVX1 INVX1_518 ( .A(cpuregs_17_[22]), .Y(_6959_) );
AOI21X1 AOI21X1_223 ( .A(decoded_rs2_0_bF_buf49_), .B(_6959_), .C(decoded_rs2_1_bF_buf10_), .Y(_6960_) );
OAI21X1 OAI21X1_992 ( .A(decoded_rs2_0_bF_buf48_), .B(cpuregs_16_[22]), .C(_6960_), .Y(_6961_) );
NOR2X1 NOR2X1_424 ( .A(cpuregs_19_[22]), .B(_5362__bF_buf14), .Y(_6962_) );
OAI21X1 OAI21X1_993 ( .A(decoded_rs2_0_bF_buf47_), .B(cpuregs_18_[22]), .C(decoded_rs2_1_bF_buf9_), .Y(_6963_) );
OAI21X1 OAI21X1_994 ( .A(_6962_), .B(_6963_), .C(_6961_), .Y(_6964_) );
INVX1 INVX1_519 ( .A(cpuregs_21_[22]), .Y(_6965_) );
AOI21X1 AOI21X1_224 ( .A(decoded_rs2_0_bF_buf46_), .B(_6965_), .C(decoded_rs2_1_bF_buf8_), .Y(_6966_) );
OAI21X1 OAI21X1_995 ( .A(decoded_rs2_0_bF_buf45_), .B(cpuregs_20_[22]), .C(_6966_), .Y(_6967_) );
INVX1 INVX1_520 ( .A(cpuregs_22_[22]), .Y(_6968_) );
AOI21X1 AOI21X1_225 ( .A(_5362__bF_buf13), .B(_6968_), .C(_5349__bF_buf11), .Y(_6969_) );
OAI21X1 OAI21X1_996 ( .A(_5362__bF_buf12), .B(cpuregs_23_[22]), .C(_6969_), .Y(_6970_) );
NAND3X1 NAND3X1_29 ( .A(decoded_rs2_2_bF_buf3_), .B(_6967_), .C(_6970_), .Y(_6971_) );
OAI21X1 OAI21X1_997 ( .A(_6964_), .B(decoded_rs2_2_bF_buf2_), .C(_6971_), .Y(_6972_) );
OAI21X1 OAI21X1_998 ( .A(decoded_rs2_3_bF_buf0_), .B(_6972_), .C(_6958_), .Y(_6973_) );
NOR2X1 NOR2X1_425 ( .A(_5347_), .B(_6973_), .Y(_6974_) );
NOR2X1 NOR2X1_426 ( .A(_5890__bF_buf3), .B(_6974_), .Y(_6975_) );
OAI21X1 OAI21X1_999 ( .A(decoded_rs2_4_bF_buf2_), .B(_6941_), .C(_6975_), .Y(_6976_) );
AOI21X1 AOI21X1_226 ( .A(decoded_imm_22_), .B(_5849__bF_buf2), .C(_4540__bF_buf4), .Y(_6977_) );
AOI22X1 AOI22X1_30 ( .A(_5224_), .B(_4540__bF_buf3), .C(_6976_), .D(_6977_), .Y(_82__22_) );
INVX1 INVX1_521 ( .A(cpuregs_1_[23]), .Y(_6978_) );
AOI21X1 AOI21X1_227 ( .A(decoded_rs2_0_bF_buf44_), .B(_6978_), .C(decoded_rs2_1_bF_buf7_), .Y(_6979_) );
OAI21X1 OAI21X1_1000 ( .A(decoded_rs2_0_bF_buf43_), .B(cpuregs_0_[23]), .C(_6979_), .Y(_6980_) );
NOR2X1 NOR2X1_427 ( .A(cpuregs_3_[23]), .B(_5362__bF_buf11), .Y(_6981_) );
OAI21X1 OAI21X1_1001 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_2_[23]), .C(decoded_rs2_1_bF_buf6_), .Y(_6982_) );
OAI21X1 OAI21X1_1002 ( .A(_6981_), .B(_6982_), .C(_6980_), .Y(_6983_) );
NOR2X1 NOR2X1_428 ( .A(decoded_rs2_0_bF_buf41_), .B(cpuregs_4_[23]), .Y(_6984_) );
OAI21X1 OAI21X1_1003 ( .A(_5362__bF_buf10), .B(cpuregs_5_[23]), .C(_5349__bF_buf10), .Y(_6985_) );
INVX1 INVX1_522 ( .A(cpuregs_6_[23]), .Y(_6986_) );
AOI21X1 AOI21X1_228 ( .A(_6986_), .B(_5362__bF_buf9), .C(_5349__bF_buf9), .Y(_6987_) );
OAI21X1 OAI21X1_1004 ( .A(cpuregs_7_[23]), .B(_5362__bF_buf8), .C(_6987_), .Y(_6988_) );
OAI21X1 OAI21X1_1005 ( .A(_6984_), .B(_6985_), .C(_6988_), .Y(_6989_) );
MUX2X1 MUX2X1_116 ( .A(_6989_), .B(_6983_), .S(decoded_rs2_2_bF_buf1_), .Y(_6990_) );
INVX1 INVX1_523 ( .A(cpuregs_8_[23]), .Y(_6991_) );
OAI21X1 OAI21X1_1006 ( .A(_5362__bF_buf7), .B(cpuregs_9_[23]), .C(_5349__bF_buf8), .Y(_6992_) );
AOI21X1 AOI21X1_229 ( .A(_6991_), .B(_5362__bF_buf6), .C(_6992_), .Y(_6993_) );
INVX1 INVX1_524 ( .A(cpuregs_10_[23]), .Y(_6994_) );
NAND2X1 NAND2X1_406 ( .A(decoded_rs2_0_bF_buf40_), .B(cpuregs_11_[23]), .Y(_6995_) );
OAI21X1 OAI21X1_1007 ( .A(_6994_), .B(decoded_rs2_0_bF_buf39_), .C(_6995_), .Y(_6996_) );
AOI21X1 AOI21X1_230 ( .A(decoded_rs2_1_bF_buf5_), .B(_6996_), .C(_6993_), .Y(_6997_) );
AND2X2 AND2X2_40 ( .A(_6997_), .B(_5358__bF_buf8), .Y(_6998_) );
INVX1 INVX1_525 ( .A(cpuregs_13_[23]), .Y(_6999_) );
AOI21X1 AOI21X1_231 ( .A(decoded_rs2_0_bF_buf38_), .B(_6999_), .C(decoded_rs2_1_bF_buf4_), .Y(_7000_) );
OAI21X1 OAI21X1_1008 ( .A(decoded_rs2_0_bF_buf37_), .B(cpuregs_12_[23]), .C(_7000_), .Y(_7001_) );
NOR2X1 NOR2X1_429 ( .A(cpuregs_15_[23]), .B(_5362__bF_buf5), .Y(_7002_) );
OAI21X1 OAI21X1_1009 ( .A(decoded_rs2_0_bF_buf36_), .B(cpuregs_14_[23]), .C(decoded_rs2_1_bF_buf3_), .Y(_7003_) );
OAI21X1 OAI21X1_1010 ( .A(_7002_), .B(_7003_), .C(_7001_), .Y(_7004_) );
OAI21X1 OAI21X1_1011 ( .A(_7004_), .B(_5358__bF_buf7), .C(decoded_rs2_3_bF_buf6_), .Y(_7005_) );
OAI22X1 OAI22X1_67 ( .A(decoded_rs2_3_bF_buf5_), .B(_6990_), .C(_6998_), .D(_7005_), .Y(_7006_) );
INVX1 INVX1_526 ( .A(cpuregs_16_[23]), .Y(_7007_) );
NAND2X1 NAND2X1_407 ( .A(decoded_rs2_0_bF_buf35_), .B(cpuregs_17_[23]), .Y(_7008_) );
OAI21X1 OAI21X1_1012 ( .A(_7007_), .B(decoded_rs2_0_bF_buf34_), .C(_7008_), .Y(_7009_) );
INVX1 INVX1_527 ( .A(cpuregs_18_[23]), .Y(_7010_) );
NAND2X1 NAND2X1_408 ( .A(decoded_rs2_0_bF_buf33_), .B(cpuregs_19_[23]), .Y(_7011_) );
OAI21X1 OAI21X1_1013 ( .A(_7010_), .B(decoded_rs2_0_bF_buf32_), .C(_7011_), .Y(_7012_) );
MUX2X1 MUX2X1_117 ( .A(_7012_), .B(_7009_), .S(decoded_rs2_1_bF_buf2_), .Y(_7013_) );
INVX1 INVX1_528 ( .A(cpuregs_20_[23]), .Y(_7014_) );
NAND2X1 NAND2X1_409 ( .A(decoded_rs2_0_bF_buf31_), .B(cpuregs_21_[23]), .Y(_7015_) );
OAI21X1 OAI21X1_1014 ( .A(_7014_), .B(decoded_rs2_0_bF_buf30_), .C(_7015_), .Y(_7016_) );
INVX1 INVX1_529 ( .A(cpuregs_22_[23]), .Y(_7017_) );
NAND2X1 NAND2X1_410 ( .A(decoded_rs2_0_bF_buf29_), .B(cpuregs_23_[23]), .Y(_7018_) );
OAI21X1 OAI21X1_1015 ( .A(_7017_), .B(decoded_rs2_0_bF_buf28_), .C(_7018_), .Y(_7019_) );
MUX2X1 MUX2X1_118 ( .A(_7019_), .B(_7016_), .S(decoded_rs2_1_bF_buf1_), .Y(_7020_) );
MUX2X1 MUX2X1_119 ( .A(_7020_), .B(_7013_), .S(decoded_rs2_2_bF_buf0_), .Y(_7021_) );
INVX1 INVX1_530 ( .A(cpuregs_28_[23]), .Y(_7022_) );
NAND2X1 NAND2X1_411 ( .A(decoded_rs2_0_bF_buf27_), .B(cpuregs_29_[23]), .Y(_7023_) );
OAI21X1 OAI21X1_1016 ( .A(_7022_), .B(decoded_rs2_0_bF_buf26_), .C(_7023_), .Y(_7024_) );
INVX1 INVX1_531 ( .A(cpuregs_31_[23]), .Y(_7025_) );
NAND2X1 NAND2X1_412 ( .A(cpuregs_30_[23]), .B(_5362__bF_buf4), .Y(_7026_) );
OAI21X1 OAI21X1_1017 ( .A(_5362__bF_buf3), .B(_7025_), .C(_7026_), .Y(_7027_) );
MUX2X1 MUX2X1_120 ( .A(_7027_), .B(_7024_), .S(decoded_rs2_1_bF_buf0_), .Y(_7028_) );
NAND2X1 NAND2X1_413 ( .A(decoded_rs2_2_bF_buf8_), .B(_7028_), .Y(_7029_) );
INVX1 INVX1_532 ( .A(cpuregs_24_[23]), .Y(_7030_) );
NAND2X1 NAND2X1_414 ( .A(decoded_rs2_0_bF_buf25_), .B(cpuregs_25_[23]), .Y(_7031_) );
OAI21X1 OAI21X1_1018 ( .A(_7030_), .B(decoded_rs2_0_bF_buf24_), .C(_7031_), .Y(_7032_) );
INVX1 INVX1_533 ( .A(cpuregs_27_[23]), .Y(_7033_) );
OAI21X1 OAI21X1_1019 ( .A(decoded_rs2_0_bF_buf23_), .B(cpuregs_26_[23]), .C(decoded_rs2_1_bF_buf45_), .Y(_7034_) );
AOI21X1 AOI21X1_232 ( .A(decoded_rs2_0_bF_buf22_), .B(_7033_), .C(_7034_), .Y(_7035_) );
AOI21X1 AOI21X1_233 ( .A(_5349__bF_buf7), .B(_7032_), .C(_7035_), .Y(_7036_) );
AOI21X1 AOI21X1_234 ( .A(_5358__bF_buf6), .B(_7036_), .C(_5348__bF_buf0), .Y(_7037_) );
AOI22X1 AOI22X1_31 ( .A(_5348__bF_buf5), .B(_7021_), .C(_7029_), .D(_7037_), .Y(_7038_) );
AOI21X1 AOI21X1_235 ( .A(decoded_rs2_4_bF_buf1_), .B(_7038_), .C(_5890__bF_buf2), .Y(_7039_) );
OAI21X1 OAI21X1_1020 ( .A(_7006_), .B(decoded_rs2_4_bF_buf0_), .C(_7039_), .Y(_7040_) );
AOI21X1 AOI21X1_236 ( .A(decoded_imm_23_), .B(_5849__bF_buf1), .C(_4540__bF_buf2), .Y(_7041_) );
AOI22X1 AOI22X1_32 ( .A(_5223_), .B(_4540__bF_buf1), .C(_7040_), .D(_7041_), .Y(_82__23_) );
INVX1 INVX1_534 ( .A(cpuregs_1_[24]), .Y(_7042_) );
AOI21X1 AOI21X1_237 ( .A(decoded_rs2_0_bF_buf21_), .B(_7042_), .C(decoded_rs2_1_bF_buf44_), .Y(_7043_) );
OAI21X1 OAI21X1_1021 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_0_[24]), .C(_7043_), .Y(_7044_) );
NOR2X1 NOR2X1_430 ( .A(cpuregs_3_[24]), .B(_5362__bF_buf2), .Y(_7045_) );
OAI21X1 OAI21X1_1022 ( .A(decoded_rs2_0_bF_buf19_), .B(cpuregs_2_[24]), .C(decoded_rs2_1_bF_buf43_), .Y(_7046_) );
OAI21X1 OAI21X1_1023 ( .A(_7045_), .B(_7046_), .C(_7044_), .Y(_7047_) );
NOR2X1 NOR2X1_431 ( .A(decoded_rs2_2_bF_buf7_), .B(_7047_), .Y(_7048_) );
INVX1 INVX1_535 ( .A(cpuregs_6_[24]), .Y(_7049_) );
AOI21X1 AOI21X1_238 ( .A(decoded_rs2_1_bF_buf42_), .B(_7049_), .C(decoded_rs2_0_bF_buf18_), .Y(_7050_) );
OAI21X1 OAI21X1_1024 ( .A(decoded_rs2_1_bF_buf41_), .B(cpuregs_4_[24]), .C(_7050_), .Y(_7051_) );
NOR2X1 NOR2X1_432 ( .A(cpuregs_5_[24]), .B(decoded_rs2_1_bF_buf40_), .Y(_7052_) );
OAI21X1 OAI21X1_1025 ( .A(_5349__bF_buf6), .B(cpuregs_7_[24]), .C(decoded_rs2_0_bF_buf17_), .Y(_7053_) );
OAI21X1 OAI21X1_1026 ( .A(_7052_), .B(_7053_), .C(_7051_), .Y(_7054_) );
OAI21X1 OAI21X1_1027 ( .A(_7054_), .B(_5358__bF_buf5), .C(_5348__bF_buf4), .Y(_7055_) );
NOR2X1 NOR2X1_433 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_12_[24]), .Y(_7056_) );
OAI21X1 OAI21X1_1028 ( .A(_5362__bF_buf1), .B(cpuregs_13_[24]), .C(_5349__bF_buf5), .Y(_7057_) );
NOR2X1 NOR2X1_434 ( .A(cpuregs_15_[24]), .B(_5362__bF_buf0), .Y(_7058_) );
OAI21X1 OAI21X1_1029 ( .A(decoded_rs2_0_bF_buf15_), .B(cpuregs_14_[24]), .C(decoded_rs2_1_bF_buf39_), .Y(_7059_) );
OAI22X1 OAI22X1_68 ( .A(_7058_), .B(_7059_), .C(_7057_), .D(_7056_), .Y(_7060_) );
NOR2X1 NOR2X1_435 ( .A(_5358__bF_buf4), .B(_7060_), .Y(_7061_) );
INVX1 INVX1_536 ( .A(cpuregs_9_[24]), .Y(_7062_) );
AOI21X1 AOI21X1_239 ( .A(decoded_rs2_0_bF_buf14_), .B(_7062_), .C(decoded_rs2_1_bF_buf38_), .Y(_7063_) );
OAI21X1 OAI21X1_1030 ( .A(cpuregs_8_[24]), .B(decoded_rs2_0_bF_buf13_), .C(_7063_), .Y(_7064_) );
NOR2X1 NOR2X1_436 ( .A(cpuregs_11_[24]), .B(_5362__bF_buf14), .Y(_7065_) );
OAI21X1 OAI21X1_1031 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_10_[24]), .C(decoded_rs2_1_bF_buf37_), .Y(_7066_) );
OAI21X1 OAI21X1_1032 ( .A(_7065_), .B(_7066_), .C(_7064_), .Y(_7067_) );
OAI21X1 OAI21X1_1033 ( .A(_7067_), .B(decoded_rs2_2_bF_buf6_), .C(decoded_rs2_3_bF_buf4_), .Y(_7068_) );
OAI22X1 OAI22X1_69 ( .A(_7055_), .B(_7048_), .C(_7061_), .D(_7068_), .Y(_7069_) );
INVX1 INVX1_537 ( .A(cpuregs_16_[24]), .Y(_7070_) );
NAND2X1 NAND2X1_415 ( .A(decoded_rs2_0_bF_buf11_), .B(cpuregs_17_[24]), .Y(_7071_) );
OAI21X1 OAI21X1_1034 ( .A(_7070_), .B(decoded_rs2_0_bF_buf10_), .C(_7071_), .Y(_7072_) );
INVX1 INVX1_538 ( .A(cpuregs_18_[24]), .Y(_7073_) );
NAND2X1 NAND2X1_416 ( .A(decoded_rs2_0_bF_buf9_), .B(cpuregs_19_[24]), .Y(_7074_) );
OAI21X1 OAI21X1_1035 ( .A(_7073_), .B(decoded_rs2_0_bF_buf8_), .C(_7074_), .Y(_7075_) );
MUX2X1 MUX2X1_121 ( .A(_7075_), .B(_7072_), .S(decoded_rs2_1_bF_buf36_), .Y(_7076_) );
INVX1 INVX1_539 ( .A(cpuregs_20_[24]), .Y(_7077_) );
NAND2X1 NAND2X1_417 ( .A(decoded_rs2_0_bF_buf7_), .B(cpuregs_21_[24]), .Y(_7078_) );
OAI21X1 OAI21X1_1036 ( .A(_7077_), .B(decoded_rs2_0_bF_buf6_), .C(_7078_), .Y(_7079_) );
INVX1 INVX1_540 ( .A(cpuregs_22_[24]), .Y(_7080_) );
NAND2X1 NAND2X1_418 ( .A(decoded_rs2_0_bF_buf5_), .B(cpuregs_23_[24]), .Y(_7081_) );
OAI21X1 OAI21X1_1037 ( .A(_7080_), .B(decoded_rs2_0_bF_buf4_), .C(_7081_), .Y(_7082_) );
MUX2X1 MUX2X1_122 ( .A(_7082_), .B(_7079_), .S(decoded_rs2_1_bF_buf35_), .Y(_7083_) );
MUX2X1 MUX2X1_123 ( .A(_7083_), .B(_7076_), .S(decoded_rs2_2_bF_buf5_), .Y(_7084_) );
INVX1 INVX1_541 ( .A(cpuregs_28_[24]), .Y(_7085_) );
NAND2X1 NAND2X1_419 ( .A(decoded_rs2_0_bF_buf3_), .B(cpuregs_29_[24]), .Y(_7086_) );
OAI21X1 OAI21X1_1038 ( .A(_7085_), .B(decoded_rs2_0_bF_buf2_), .C(_7086_), .Y(_7087_) );
INVX1 INVX1_542 ( .A(cpuregs_31_[24]), .Y(_7088_) );
NAND2X1 NAND2X1_420 ( .A(cpuregs_30_[24]), .B(_5362__bF_buf13), .Y(_7089_) );
OAI21X1 OAI21X1_1039 ( .A(_5362__bF_buf12), .B(_7088_), .C(_7089_), .Y(_7090_) );
MUX2X1 MUX2X1_124 ( .A(_7090_), .B(_7087_), .S(decoded_rs2_1_bF_buf34_), .Y(_7091_) );
NAND2X1 NAND2X1_421 ( .A(decoded_rs2_2_bF_buf4_), .B(_7091_), .Y(_7092_) );
INVX1 INVX1_543 ( .A(cpuregs_24_[24]), .Y(_7093_) );
NAND2X1 NAND2X1_422 ( .A(decoded_rs2_0_bF_buf1_), .B(cpuregs_25_[24]), .Y(_7094_) );
OAI21X1 OAI21X1_1040 ( .A(_7093_), .B(decoded_rs2_0_bF_buf0_), .C(_7094_), .Y(_7095_) );
INVX1 INVX1_544 ( .A(cpuregs_27_[24]), .Y(_7096_) );
OAI21X1 OAI21X1_1041 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_26_[24]), .C(decoded_rs2_1_bF_buf33_), .Y(_7097_) );
AOI21X1 AOI21X1_240 ( .A(decoded_rs2_0_bF_buf77_), .B(_7096_), .C(_7097_), .Y(_7098_) );
AOI21X1 AOI21X1_241 ( .A(_5349__bF_buf4), .B(_7095_), .C(_7098_), .Y(_7099_) );
AOI21X1 AOI21X1_242 ( .A(_5358__bF_buf3), .B(_7099_), .C(_5348__bF_buf3), .Y(_7100_) );
AOI22X1 AOI22X1_33 ( .A(_5348__bF_buf2), .B(_7084_), .C(_7092_), .D(_7100_), .Y(_7101_) );
AOI21X1 AOI21X1_243 ( .A(decoded_rs2_4_bF_buf7_), .B(_7101_), .C(_5890__bF_buf1), .Y(_7102_) );
OAI21X1 OAI21X1_1042 ( .A(decoded_rs2_4_bF_buf6_), .B(_7069_), .C(_7102_), .Y(_7103_) );
AOI21X1 AOI21X1_244 ( .A(decoded_imm_24_), .B(_5849__bF_buf0), .C(_4540__bF_buf0), .Y(_7104_) );
AOI22X1 AOI22X1_34 ( .A(_5033_), .B(_4540__bF_buf6), .C(_7103_), .D(_7104_), .Y(_82__24_) );
INVX1 INVX1_545 ( .A(cpuregs_0_[25]), .Y(_7105_) );
NAND2X1 NAND2X1_423 ( .A(decoded_rs2_0_bF_buf76_), .B(cpuregs_1_[25]), .Y(_7106_) );
OAI21X1 OAI21X1_1043 ( .A(_7105_), .B(decoded_rs2_0_bF_buf75_), .C(_7106_), .Y(_7107_) );
INVX1 INVX1_546 ( .A(cpuregs_2_[25]), .Y(_7108_) );
NAND2X1 NAND2X1_424 ( .A(decoded_rs2_0_bF_buf74_), .B(cpuregs_3_[25]), .Y(_7109_) );
OAI21X1 OAI21X1_1044 ( .A(_7108_), .B(decoded_rs2_0_bF_buf73_), .C(_7109_), .Y(_7110_) );
MUX2X1 MUX2X1_125 ( .A(_7110_), .B(_7107_), .S(decoded_rs2_1_bF_buf32_), .Y(_7111_) );
NAND2X1 NAND2X1_425 ( .A(_5358__bF_buf2), .B(_7111_), .Y(_7112_) );
NOR2X1 NOR2X1_437 ( .A(decoded_rs2_0_bF_buf72_), .B(cpuregs_4_[25]), .Y(_7113_) );
OAI21X1 OAI21X1_1045 ( .A(_5362__bF_buf11), .B(cpuregs_5_[25]), .C(_5349__bF_buf3), .Y(_7114_) );
NOR2X1 NOR2X1_438 ( .A(cpuregs_7_[25]), .B(_5362__bF_buf10), .Y(_7115_) );
OAI21X1 OAI21X1_1046 ( .A(cpuregs_6_[25]), .B(decoded_rs2_0_bF_buf71_), .C(decoded_rs2_1_bF_buf31_), .Y(_7116_) );
OAI22X1 OAI22X1_70 ( .A(_7115_), .B(_7116_), .C(_7114_), .D(_7113_), .Y(_7117_) );
OAI21X1 OAI21X1_1047 ( .A(_5358__bF_buf1), .B(_7117_), .C(_7112_), .Y(_7118_) );
INVX1 INVX1_547 ( .A(cpuregs_9_[25]), .Y(_7119_) );
AOI21X1 AOI21X1_245 ( .A(decoded_rs2_0_bF_buf70_), .B(_7119_), .C(decoded_rs2_1_bF_buf30_), .Y(_7120_) );
OAI21X1 OAI21X1_1048 ( .A(cpuregs_8_[25]), .B(decoded_rs2_0_bF_buf69_), .C(_7120_), .Y(_7121_) );
NOR2X1 NOR2X1_439 ( .A(cpuregs_11_[25]), .B(_5362__bF_buf9), .Y(_7122_) );
OAI21X1 OAI21X1_1049 ( .A(decoded_rs2_0_bF_buf68_), .B(cpuregs_10_[25]), .C(decoded_rs2_1_bF_buf29_), .Y(_7123_) );
OAI21X1 OAI21X1_1050 ( .A(_7122_), .B(_7123_), .C(_7121_), .Y(_7124_) );
INVX1 INVX1_548 ( .A(cpuregs_12_[25]), .Y(_7125_) );
NAND2X1 NAND2X1_426 ( .A(decoded_rs2_0_bF_buf67_), .B(cpuregs_13_[25]), .Y(_7126_) );
OAI21X1 OAI21X1_1051 ( .A(_7125_), .B(decoded_rs2_0_bF_buf66_), .C(_7126_), .Y(_7127_) );
INVX1 INVX1_549 ( .A(cpuregs_15_[25]), .Y(_7128_) );
OAI21X1 OAI21X1_1052 ( .A(decoded_rs2_0_bF_buf65_), .B(cpuregs_14_[25]), .C(decoded_rs2_1_bF_buf28_), .Y(_7129_) );
AOI21X1 AOI21X1_246 ( .A(decoded_rs2_0_bF_buf64_), .B(_7128_), .C(_7129_), .Y(_7130_) );
AOI21X1 AOI21X1_247 ( .A(_5349__bF_buf2), .B(_7127_), .C(_7130_), .Y(_7131_) );
AOI21X1 AOI21X1_248 ( .A(decoded_rs2_2_bF_buf3_), .B(_7131_), .C(_5348__bF_buf1), .Y(_7132_) );
OAI21X1 OAI21X1_1053 ( .A(decoded_rs2_2_bF_buf2_), .B(_7124_), .C(_7132_), .Y(_7133_) );
OAI21X1 OAI21X1_1054 ( .A(_7118_), .B(decoded_rs2_3_bF_buf3_), .C(_7133_), .Y(_7134_) );
INVX1 INVX1_550 ( .A(cpuregs_26_[25]), .Y(_7135_) );
OAI21X1 OAI21X1_1055 ( .A(_7135_), .B(decoded_rs2_0_bF_buf63_), .C(decoded_rs2_1_bF_buf27_), .Y(_7136_) );
AOI21X1 AOI21X1_249 ( .A(decoded_rs2_0_bF_buf62_), .B(cpuregs_27_[25]), .C(_7136_), .Y(_7137_) );
AND2X2 AND2X2_41 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_25_[25]), .Y(_7138_) );
INVX1 INVX1_551 ( .A(cpuregs_24_[25]), .Y(_7139_) );
OAI21X1 OAI21X1_1056 ( .A(_7139_), .B(decoded_rs2_0_bF_buf60_), .C(_5349__bF_buf1), .Y(_7140_) );
OAI21X1 OAI21X1_1057 ( .A(_7140_), .B(_7138_), .C(_5358__bF_buf0), .Y(_7141_) );
INVX1 INVX1_552 ( .A(cpuregs_29_[25]), .Y(_7142_) );
NAND2X1 NAND2X1_427 ( .A(cpuregs_28_[25]), .B(_5362__bF_buf8), .Y(_7143_) );
OAI21X1 OAI21X1_1058 ( .A(_5362__bF_buf7), .B(_7142_), .C(_7143_), .Y(_7144_) );
INVX1 INVX1_553 ( .A(cpuregs_31_[25]), .Y(_7145_) );
OAI21X1 OAI21X1_1059 ( .A(decoded_rs2_0_bF_buf59_), .B(cpuregs_30_[25]), .C(decoded_rs2_1_bF_buf26_), .Y(_7146_) );
AOI21X1 AOI21X1_250 ( .A(decoded_rs2_0_bF_buf58_), .B(_7145_), .C(_7146_), .Y(_7147_) );
AOI21X1 AOI21X1_251 ( .A(_5349__bF_buf0), .B(_7144_), .C(_7147_), .Y(_7148_) );
OAI22X1 OAI22X1_71 ( .A(_7141_), .B(_7137_), .C(_7148_), .D(_5358__bF_buf12), .Y(_7149_) );
INVX1 INVX1_554 ( .A(cpuregs_16_[25]), .Y(_7150_) );
NAND2X1 NAND2X1_428 ( .A(decoded_rs2_0_bF_buf57_), .B(cpuregs_17_[25]), .Y(_7151_) );
OAI21X1 OAI21X1_1060 ( .A(_7150_), .B(decoded_rs2_0_bF_buf56_), .C(_7151_), .Y(_7152_) );
INVX1 INVX1_555 ( .A(cpuregs_19_[25]), .Y(_7153_) );
OAI21X1 OAI21X1_1061 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_18_[25]), .C(decoded_rs2_1_bF_buf25_), .Y(_7154_) );
AOI21X1 AOI21X1_252 ( .A(decoded_rs2_0_bF_buf54_), .B(_7153_), .C(_7154_), .Y(_7155_) );
AOI21X1 AOI21X1_253 ( .A(_5349__bF_buf11), .B(_7152_), .C(_7155_), .Y(_7156_) );
NAND2X1 NAND2X1_429 ( .A(_5358__bF_buf11), .B(_7156_), .Y(_7157_) );
INVX1 INVX1_556 ( .A(cpuregs_20_[25]), .Y(_7158_) );
NAND2X1 NAND2X1_430 ( .A(decoded_rs2_0_bF_buf53_), .B(cpuregs_21_[25]), .Y(_7159_) );
OAI21X1 OAI21X1_1062 ( .A(_7158_), .B(decoded_rs2_0_bF_buf52_), .C(_7159_), .Y(_7160_) );
INVX1 INVX1_557 ( .A(cpuregs_22_[25]), .Y(_7161_) );
NAND2X1 NAND2X1_431 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_23_[25]), .Y(_7162_) );
OAI21X1 OAI21X1_1063 ( .A(_7161_), .B(decoded_rs2_0_bF_buf50_), .C(_7162_), .Y(_7163_) );
MUX2X1 MUX2X1_126 ( .A(_7163_), .B(_7160_), .S(decoded_rs2_1_bF_buf24_), .Y(_7164_) );
AOI21X1 AOI21X1_254 ( .A(decoded_rs2_2_bF_buf1_), .B(_7164_), .C(decoded_rs2_3_bF_buf2_), .Y(_7165_) );
AOI22X1 AOI22X1_35 ( .A(_7165_), .B(_7157_), .C(decoded_rs2_3_bF_buf1_), .D(_7149_), .Y(_7166_) );
AOI21X1 AOI21X1_255 ( .A(decoded_rs2_4_bF_buf5_), .B(_7166_), .C(_5890__bF_buf0), .Y(_7167_) );
OAI21X1 OAI21X1_1064 ( .A(decoded_rs2_4_bF_buf4_), .B(_7134_), .C(_7167_), .Y(_7168_) );
AOI21X1 AOI21X1_256 ( .A(decoded_imm_25_), .B(_5849__bF_buf4), .C(_4540__bF_buf5), .Y(_7169_) );
AOI22X1 AOI22X1_36 ( .A(_5028_), .B(_4540__bF_buf4), .C(_7168_), .D(_7169_), .Y(_82__25_) );
INVX1 INVX1_558 ( .A(cpuregs_1_[26]), .Y(_7170_) );
AOI21X1 AOI21X1_257 ( .A(decoded_rs2_0_bF_buf49_), .B(_7170_), .C(decoded_rs2_1_bF_buf23_), .Y(_7171_) );
OAI21X1 OAI21X1_1065 ( .A(decoded_rs2_0_bF_buf48_), .B(cpuregs_0_[26]), .C(_7171_), .Y(_7172_) );
NOR2X1 NOR2X1_440 ( .A(cpuregs_3_[26]), .B(_5362__bF_buf6), .Y(_7173_) );
OAI21X1 OAI21X1_1066 ( .A(decoded_rs2_0_bF_buf47_), .B(cpuregs_2_[26]), .C(decoded_rs2_1_bF_buf22_), .Y(_7174_) );
OAI21X1 OAI21X1_1067 ( .A(_7173_), .B(_7174_), .C(_7172_), .Y(_7175_) );
NOR2X1 NOR2X1_441 ( .A(decoded_rs2_2_bF_buf0_), .B(_7175_), .Y(_7176_) );
NOR2X1 NOR2X1_442 ( .A(decoded_rs2_0_bF_buf46_), .B(cpuregs_4_[26]), .Y(_7177_) );
OAI21X1 OAI21X1_1068 ( .A(_5362__bF_buf5), .B(cpuregs_5_[26]), .C(_5349__bF_buf10), .Y(_7178_) );
NOR2X1 NOR2X1_443 ( .A(cpuregs_7_[26]), .B(_5362__bF_buf4), .Y(_7179_) );
OAI21X1 OAI21X1_1069 ( .A(cpuregs_6_[26]), .B(decoded_rs2_0_bF_buf45_), .C(decoded_rs2_1_bF_buf21_), .Y(_7180_) );
OAI22X1 OAI22X1_72 ( .A(_7179_), .B(_7180_), .C(_7178_), .D(_7177_), .Y(_7181_) );
OAI21X1 OAI21X1_1070 ( .A(_7181_), .B(_5358__bF_buf10), .C(_5348__bF_buf0), .Y(_7182_) );
INVX1 INVX1_559 ( .A(cpuregs_13_[26]), .Y(_7183_) );
AOI21X1 AOI21X1_258 ( .A(decoded_rs2_0_bF_buf44_), .B(_7183_), .C(decoded_rs2_1_bF_buf20_), .Y(_7184_) );
OAI21X1 OAI21X1_1071 ( .A(decoded_rs2_0_bF_buf43_), .B(cpuregs_12_[26]), .C(_7184_), .Y(_7185_) );
NOR2X1 NOR2X1_444 ( .A(cpuregs_15_[26]), .B(_5362__bF_buf3), .Y(_7186_) );
OAI21X1 OAI21X1_1072 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_14_[26]), .C(decoded_rs2_1_bF_buf19_), .Y(_7187_) );
OAI21X1 OAI21X1_1073 ( .A(_7186_), .B(_7187_), .C(_7185_), .Y(_7188_) );
NOR2X1 NOR2X1_445 ( .A(_5358__bF_buf9), .B(_7188_), .Y(_7189_) );
NOR2X1 NOR2X1_446 ( .A(cpuregs_8_[26]), .B(decoded_rs2_0_bF_buf41_), .Y(_7190_) );
OAI21X1 OAI21X1_1074 ( .A(_5362__bF_buf2), .B(cpuregs_9_[26]), .C(_5349__bF_buf9), .Y(_7191_) );
NOR2X1 NOR2X1_447 ( .A(cpuregs_11_[26]), .B(_5362__bF_buf1), .Y(_7192_) );
OAI21X1 OAI21X1_1075 ( .A(decoded_rs2_0_bF_buf40_), .B(cpuregs_10_[26]), .C(decoded_rs2_1_bF_buf18_), .Y(_7193_) );
OAI22X1 OAI22X1_73 ( .A(_7192_), .B(_7193_), .C(_7191_), .D(_7190_), .Y(_7194_) );
OAI21X1 OAI21X1_1076 ( .A(_7194_), .B(decoded_rs2_2_bF_buf8_), .C(decoded_rs2_3_bF_buf0_), .Y(_7195_) );
OAI22X1 OAI22X1_74 ( .A(_7176_), .B(_7182_), .C(_7195_), .D(_7189_), .Y(_7196_) );
INVX1 INVX1_560 ( .A(cpuregs_26_[26]), .Y(_7197_) );
OAI21X1 OAI21X1_1077 ( .A(_7197_), .B(decoded_rs2_0_bF_buf39_), .C(decoded_rs2_1_bF_buf17_), .Y(_7198_) );
AOI21X1 AOI21X1_259 ( .A(decoded_rs2_0_bF_buf38_), .B(cpuregs_27_[26]), .C(_7198_), .Y(_7199_) );
AND2X2 AND2X2_42 ( .A(decoded_rs2_0_bF_buf37_), .B(cpuregs_25_[26]), .Y(_7200_) );
INVX1 INVX1_561 ( .A(cpuregs_24_[26]), .Y(_7201_) );
OAI21X1 OAI21X1_1078 ( .A(_7201_), .B(decoded_rs2_0_bF_buf36_), .C(_5349__bF_buf8), .Y(_7202_) );
OAI21X1 OAI21X1_1079 ( .A(_7202_), .B(_7200_), .C(_5358__bF_buf8), .Y(_7203_) );
INVX1 INVX1_562 ( .A(cpuregs_30_[26]), .Y(_7204_) );
OAI21X1 OAI21X1_1080 ( .A(_7204_), .B(decoded_rs2_0_bF_buf35_), .C(decoded_rs2_1_bF_buf16_), .Y(_7205_) );
AOI21X1 AOI21X1_260 ( .A(decoded_rs2_0_bF_buf34_), .B(cpuregs_31_[26]), .C(_7205_), .Y(_7206_) );
INVX1 INVX1_563 ( .A(cpuregs_28_[26]), .Y(_7207_) );
NOR2X1 NOR2X1_448 ( .A(decoded_rs2_0_bF_buf33_), .B(_7207_), .Y(_7208_) );
INVX1 INVX1_564 ( .A(cpuregs_29_[26]), .Y(_7209_) );
OAI21X1 OAI21X1_1081 ( .A(_5362__bF_buf0), .B(_7209_), .C(_5349__bF_buf7), .Y(_7210_) );
OAI21X1 OAI21X1_1082 ( .A(_7210_), .B(_7208_), .C(decoded_rs2_2_bF_buf7_), .Y(_7211_) );
OAI22X1 OAI22X1_75 ( .A(_7203_), .B(_7199_), .C(_7211_), .D(_7206_), .Y(_7212_) );
INVX1 INVX1_565 ( .A(cpuregs_17_[26]), .Y(_7213_) );
NAND2X1 NAND2X1_432 ( .A(cpuregs_16_[26]), .B(_5362__bF_buf14), .Y(_7214_) );
OAI21X1 OAI21X1_1083 ( .A(_5362__bF_buf13), .B(_7213_), .C(_7214_), .Y(_7215_) );
INVX1 INVX1_566 ( .A(cpuregs_19_[26]), .Y(_7216_) );
OAI21X1 OAI21X1_1084 ( .A(decoded_rs2_0_bF_buf32_), .B(cpuregs_18_[26]), .C(decoded_rs2_1_bF_buf15_), .Y(_7217_) );
AOI21X1 AOI21X1_261 ( .A(decoded_rs2_0_bF_buf31_), .B(_7216_), .C(_7217_), .Y(_7218_) );
AOI21X1 AOI21X1_262 ( .A(_5349__bF_buf6), .B(_7215_), .C(_7218_), .Y(_7219_) );
NAND2X1 NAND2X1_433 ( .A(_5358__bF_buf7), .B(_7219_), .Y(_7220_) );
INVX1 INVX1_567 ( .A(cpuregs_20_[26]), .Y(_7221_) );
NAND2X1 NAND2X1_434 ( .A(decoded_rs2_0_bF_buf30_), .B(cpuregs_21_[26]), .Y(_7222_) );
OAI21X1 OAI21X1_1085 ( .A(_7221_), .B(decoded_rs2_0_bF_buf29_), .C(_7222_), .Y(_7223_) );
INVX1 INVX1_568 ( .A(cpuregs_22_[26]), .Y(_7224_) );
NAND2X1 NAND2X1_435 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_23_[26]), .Y(_7225_) );
OAI21X1 OAI21X1_1086 ( .A(_7224_), .B(decoded_rs2_0_bF_buf27_), .C(_7225_), .Y(_7226_) );
MUX2X1 MUX2X1_127 ( .A(_7226_), .B(_7223_), .S(decoded_rs2_1_bF_buf14_), .Y(_7227_) );
AOI21X1 AOI21X1_263 ( .A(decoded_rs2_2_bF_buf6_), .B(_7227_), .C(decoded_rs2_3_bF_buf6_), .Y(_7228_) );
AOI22X1 AOI22X1_37 ( .A(_7228_), .B(_7220_), .C(decoded_rs2_3_bF_buf5_), .D(_7212_), .Y(_7229_) );
AOI21X1 AOI21X1_264 ( .A(decoded_rs2_4_bF_buf3_), .B(_7229_), .C(_5890__bF_buf3), .Y(_7230_) );
OAI21X1 OAI21X1_1087 ( .A(decoded_rs2_4_bF_buf2_), .B(_7196_), .C(_7230_), .Y(_7231_) );
AOI21X1 AOI21X1_265 ( .A(decoded_imm_26_), .B(_5849__bF_buf3), .C(_4540__bF_buf3), .Y(_7232_) );
AOI22X1 AOI22X1_38 ( .A(_5022_), .B(_4540__bF_buf2), .C(_7231_), .D(_7232_), .Y(_82__26_) );
INVX1 INVX1_569 ( .A(cpuregs_2_[27]), .Y(_7233_) );
AOI21X1 AOI21X1_266 ( .A(decoded_rs2_1_bF_buf13_), .B(_7233_), .C(decoded_rs2_0_bF_buf26_), .Y(_7234_) );
OAI21X1 OAI21X1_1088 ( .A(decoded_rs2_1_bF_buf12_), .B(cpuregs_0_[27]), .C(_7234_), .Y(_7235_) );
NOR2X1 NOR2X1_449 ( .A(decoded_rs2_1_bF_buf11_), .B(cpuregs_1_[27]), .Y(_7236_) );
OAI21X1 OAI21X1_1089 ( .A(_5349__bF_buf5), .B(cpuregs_3_[27]), .C(decoded_rs2_0_bF_buf25_), .Y(_7237_) );
OAI21X1 OAI21X1_1090 ( .A(_7236_), .B(_7237_), .C(_7235_), .Y(_7238_) );
NOR2X1 NOR2X1_450 ( .A(decoded_rs2_2_bF_buf5_), .B(_7238_), .Y(_7239_) );
INVX1 INVX1_570 ( .A(cpuregs_6_[27]), .Y(_7240_) );
AOI21X1 AOI21X1_267 ( .A(decoded_rs2_1_bF_buf10_), .B(_7240_), .C(decoded_rs2_0_bF_buf24_), .Y(_7241_) );
OAI21X1 OAI21X1_1091 ( .A(decoded_rs2_1_bF_buf9_), .B(cpuregs_4_[27]), .C(_7241_), .Y(_7242_) );
NOR2X1 NOR2X1_451 ( .A(cpuregs_5_[27]), .B(decoded_rs2_1_bF_buf8_), .Y(_7243_) );
OAI21X1 OAI21X1_1092 ( .A(_5349__bF_buf4), .B(cpuregs_7_[27]), .C(decoded_rs2_0_bF_buf23_), .Y(_7244_) );
OAI21X1 OAI21X1_1093 ( .A(_7243_), .B(_7244_), .C(_7242_), .Y(_7245_) );
OAI21X1 OAI21X1_1094 ( .A(_7245_), .B(_5358__bF_buf6), .C(_5348__bF_buf5), .Y(_7246_) );
INVX1 INVX1_571 ( .A(cpuregs_13_[27]), .Y(_7247_) );
AOI21X1 AOI21X1_268 ( .A(decoded_rs2_0_bF_buf22_), .B(_7247_), .C(decoded_rs2_1_bF_buf7_), .Y(_7248_) );
OAI21X1 OAI21X1_1095 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_12_[27]), .C(_7248_), .Y(_7249_) );
NOR2X1 NOR2X1_452 ( .A(cpuregs_15_[27]), .B(_5362__bF_buf12), .Y(_7250_) );
OAI21X1 OAI21X1_1096 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_14_[27]), .C(decoded_rs2_1_bF_buf6_), .Y(_7251_) );
OAI21X1 OAI21X1_1097 ( .A(_7250_), .B(_7251_), .C(_7249_), .Y(_7252_) );
NOR2X1 NOR2X1_453 ( .A(_5358__bF_buf5), .B(_7252_), .Y(_7253_) );
INVX1 INVX1_572 ( .A(cpuregs_9_[27]), .Y(_7254_) );
AOI21X1 AOI21X1_269 ( .A(decoded_rs2_0_bF_buf19_), .B(_7254_), .C(decoded_rs2_1_bF_buf5_), .Y(_7255_) );
OAI21X1 OAI21X1_1098 ( .A(cpuregs_8_[27]), .B(decoded_rs2_0_bF_buf18_), .C(_7255_), .Y(_7256_) );
NOR2X1 NOR2X1_454 ( .A(cpuregs_11_[27]), .B(_5362__bF_buf11), .Y(_7257_) );
OAI21X1 OAI21X1_1099 ( .A(decoded_rs2_0_bF_buf17_), .B(cpuregs_10_[27]), .C(decoded_rs2_1_bF_buf4_), .Y(_7258_) );
OAI21X1 OAI21X1_1100 ( .A(_7257_), .B(_7258_), .C(_7256_), .Y(_7259_) );
OAI21X1 OAI21X1_1101 ( .A(_7259_), .B(decoded_rs2_2_bF_buf4_), .C(decoded_rs2_3_bF_buf4_), .Y(_7260_) );
OAI22X1 OAI22X1_76 ( .A(_7246_), .B(_7239_), .C(_7253_), .D(_7260_), .Y(_7261_) );
INVX1 INVX1_573 ( .A(cpuregs_26_[27]), .Y(_7262_) );
OAI21X1 OAI21X1_1102 ( .A(_7262_), .B(decoded_rs2_0_bF_buf16_), .C(decoded_rs2_1_bF_buf3_), .Y(_7263_) );
AOI21X1 AOI21X1_270 ( .A(decoded_rs2_0_bF_buf15_), .B(cpuregs_27_[27]), .C(_7263_), .Y(_7264_) );
AND2X2 AND2X2_43 ( .A(decoded_rs2_0_bF_buf14_), .B(cpuregs_25_[27]), .Y(_7265_) );
INVX1 INVX1_574 ( .A(cpuregs_24_[27]), .Y(_7266_) );
OAI21X1 OAI21X1_1103 ( .A(_7266_), .B(decoded_rs2_0_bF_buf13_), .C(_5349__bF_buf3), .Y(_7267_) );
OAI21X1 OAI21X1_1104 ( .A(_7267_), .B(_7265_), .C(_5358__bF_buf4), .Y(_7268_) );
INVX1 INVX1_575 ( .A(cpuregs_28_[27]), .Y(_7269_) );
NAND2X1 NAND2X1_436 ( .A(decoded_rs2_0_bF_buf12_), .B(cpuregs_29_[27]), .Y(_7270_) );
OAI21X1 OAI21X1_1105 ( .A(_7269_), .B(decoded_rs2_0_bF_buf11_), .C(_7270_), .Y(_7271_) );
INVX1 INVX1_576 ( .A(cpuregs_30_[27]), .Y(_7272_) );
NAND2X1 NAND2X1_437 ( .A(decoded_rs2_0_bF_buf10_), .B(cpuregs_31_[27]), .Y(_7273_) );
OAI21X1 OAI21X1_1106 ( .A(_7272_), .B(decoded_rs2_0_bF_buf9_), .C(_7273_), .Y(_7274_) );
MUX2X1 MUX2X1_128 ( .A(_7274_), .B(_7271_), .S(decoded_rs2_1_bF_buf2_), .Y(_7275_) );
OAI22X1 OAI22X1_77 ( .A(_7268_), .B(_7264_), .C(_7275_), .D(_5358__bF_buf3), .Y(_7276_) );
INVX1 INVX1_577 ( .A(cpuregs_16_[27]), .Y(_7277_) );
NAND2X1 NAND2X1_438 ( .A(decoded_rs2_0_bF_buf8_), .B(cpuregs_17_[27]), .Y(_7278_) );
OAI21X1 OAI21X1_1107 ( .A(_7277_), .B(decoded_rs2_0_bF_buf7_), .C(_7278_), .Y(_7279_) );
INVX1 INVX1_578 ( .A(cpuregs_19_[27]), .Y(_7280_) );
OAI21X1 OAI21X1_1108 ( .A(decoded_rs2_0_bF_buf6_), .B(cpuregs_18_[27]), .C(decoded_rs2_1_bF_buf1_), .Y(_7281_) );
AOI21X1 AOI21X1_271 ( .A(decoded_rs2_0_bF_buf5_), .B(_7280_), .C(_7281_), .Y(_7282_) );
AOI21X1 AOI21X1_272 ( .A(_5349__bF_buf2), .B(_7279_), .C(_7282_), .Y(_7283_) );
NAND2X1 NAND2X1_439 ( .A(_5358__bF_buf2), .B(_7283_), .Y(_7284_) );
INVX1 INVX1_579 ( .A(cpuregs_20_[27]), .Y(_7285_) );
NAND2X1 NAND2X1_440 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_21_[27]), .Y(_7286_) );
OAI21X1 OAI21X1_1109 ( .A(_7285_), .B(decoded_rs2_0_bF_buf3_), .C(_7286_), .Y(_7287_) );
INVX1 INVX1_580 ( .A(cpuregs_22_[27]), .Y(_7288_) );
NAND2X1 NAND2X1_441 ( .A(decoded_rs2_0_bF_buf2_), .B(cpuregs_23_[27]), .Y(_7289_) );
OAI21X1 OAI21X1_1110 ( .A(_7288_), .B(decoded_rs2_0_bF_buf1_), .C(_7289_), .Y(_7290_) );
MUX2X1 MUX2X1_129 ( .A(_7290_), .B(_7287_), .S(decoded_rs2_1_bF_buf0_), .Y(_7291_) );
AOI21X1 AOI21X1_273 ( .A(decoded_rs2_2_bF_buf3_), .B(_7291_), .C(decoded_rs2_3_bF_buf3_), .Y(_7292_) );
AOI22X1 AOI22X1_39 ( .A(_7292_), .B(_7284_), .C(decoded_rs2_3_bF_buf2_), .D(_7276_), .Y(_7293_) );
AOI21X1 AOI21X1_274 ( .A(decoded_rs2_4_bF_buf1_), .B(_7293_), .C(_5890__bF_buf2), .Y(_7294_) );
OAI21X1 OAI21X1_1111 ( .A(decoded_rs2_4_bF_buf0_), .B(_7261_), .C(_7294_), .Y(_7295_) );
AOI21X1 AOI21X1_275 ( .A(decoded_imm_27_), .B(_5849__bF_buf2), .C(_4540__bF_buf1), .Y(_7296_) );
AOI22X1 AOI22X1_40 ( .A(_5017_), .B(_4540__bF_buf0), .C(_7295_), .D(_7296_), .Y(_82__27_) );
INVX1 INVX1_581 ( .A(cpuregs_20_[28]), .Y(_7297_) );
OAI21X1 OAI21X1_1112 ( .A(_5358__bF_buf1), .B(_7297_), .C(_5362__bF_buf10), .Y(_7298_) );
AOI21X1 AOI21X1_276 ( .A(_5358__bF_buf0), .B(cpuregs_16_[28]), .C(_7298_), .Y(_7299_) );
INVX1 INVX1_582 ( .A(cpuregs_21_[28]), .Y(_7300_) );
OAI21X1 OAI21X1_1113 ( .A(_5358__bF_buf12), .B(_7300_), .C(decoded_rs2_0_bF_buf0_), .Y(_7301_) );
AOI21X1 AOI21X1_277 ( .A(_5358__bF_buf11), .B(cpuregs_17_[28]), .C(_7301_), .Y(_7302_) );
OAI21X1 OAI21X1_1114 ( .A(_7299_), .B(_7302_), .C(_5349__bF_buf1), .Y(_7303_) );
INVX1 INVX1_583 ( .A(cpuregs_22_[28]), .Y(_7304_) );
OAI21X1 OAI21X1_1115 ( .A(_5358__bF_buf10), .B(_7304_), .C(_5362__bF_buf9), .Y(_7305_) );
AOI21X1 AOI21X1_278 ( .A(_5358__bF_buf9), .B(cpuregs_18_[28]), .C(_7305_), .Y(_7306_) );
INVX1 INVX1_584 ( .A(cpuregs_23_[28]), .Y(_7307_) );
OAI21X1 OAI21X1_1116 ( .A(_5358__bF_buf8), .B(_7307_), .C(decoded_rs2_0_bF_buf78_), .Y(_7308_) );
AOI21X1 AOI21X1_279 ( .A(_5358__bF_buf7), .B(cpuregs_19_[28]), .C(_7308_), .Y(_7309_) );
OAI21X1 OAI21X1_1117 ( .A(_7306_), .B(_7309_), .C(decoded_rs2_1_bF_buf45_), .Y(_7310_) );
NAND3X1 NAND3X1_30 ( .A(decoded_rs2_4_bF_buf7_), .B(_7303_), .C(_7310_), .Y(_7311_) );
INVX1 INVX1_585 ( .A(cpuregs_6_[28]), .Y(_7312_) );
AOI21X1 AOI21X1_280 ( .A(decoded_rs2_1_bF_buf44_), .B(_7312_), .C(decoded_rs2_0_bF_buf77_), .Y(_7313_) );
OAI21X1 OAI21X1_1118 ( .A(decoded_rs2_1_bF_buf43_), .B(cpuregs_4_[28]), .C(_7313_), .Y(_7314_) );
NOR2X1 NOR2X1_455 ( .A(cpuregs_5_[28]), .B(decoded_rs2_1_bF_buf42_), .Y(_7315_) );
OAI21X1 OAI21X1_1119 ( .A(_5349__bF_buf0), .B(cpuregs_7_[28]), .C(decoded_rs2_0_bF_buf76_), .Y(_7316_) );
OAI21X1 OAI21X1_1120 ( .A(_7315_), .B(_7316_), .C(_7314_), .Y(_7317_) );
INVX1 INVX1_586 ( .A(cpuregs_2_[28]), .Y(_7318_) );
AOI21X1 AOI21X1_281 ( .A(decoded_rs2_1_bF_buf41_), .B(_7318_), .C(decoded_rs2_0_bF_buf75_), .Y(_7319_) );
OAI21X1 OAI21X1_1121 ( .A(decoded_rs2_1_bF_buf40_), .B(cpuregs_0_[28]), .C(_7319_), .Y(_7320_) );
NOR2X1 NOR2X1_456 ( .A(decoded_rs2_1_bF_buf39_), .B(cpuregs_1_[28]), .Y(_7321_) );
OAI21X1 OAI21X1_1122 ( .A(_5349__bF_buf11), .B(cpuregs_3_[28]), .C(decoded_rs2_0_bF_buf74_), .Y(_7322_) );
OAI21X1 OAI21X1_1123 ( .A(_7321_), .B(_7322_), .C(_7320_), .Y(_7323_) );
MUX2X1 MUX2X1_130 ( .A(_7323_), .B(_7317_), .S(_5358__bF_buf6), .Y(_7324_) );
OAI21X1 OAI21X1_1124 ( .A(decoded_rs2_4_bF_buf6_), .B(_7324_), .C(_7311_), .Y(_7325_) );
AND2X2 AND2X2_44 ( .A(_7325_), .B(_5348__bF_buf4), .Y(_7326_) );
INVX1 INVX1_587 ( .A(cpuregs_28_[28]), .Y(_7327_) );
NAND2X1 NAND2X1_442 ( .A(decoded_rs2_0_bF_buf73_), .B(cpuregs_29_[28]), .Y(_7328_) );
OAI21X1 OAI21X1_1125 ( .A(_7327_), .B(decoded_rs2_0_bF_buf72_), .C(_7328_), .Y(_7329_) );
INVX1 INVX1_588 ( .A(cpuregs_31_[28]), .Y(_7330_) );
OAI21X1 OAI21X1_1126 ( .A(decoded_rs2_0_bF_buf71_), .B(cpuregs_30_[28]), .C(decoded_rs2_1_bF_buf38_), .Y(_7331_) );
AOI21X1 AOI21X1_282 ( .A(decoded_rs2_0_bF_buf70_), .B(_7330_), .C(_7331_), .Y(_7332_) );
AOI21X1 AOI21X1_283 ( .A(_5349__bF_buf10), .B(_7329_), .C(_7332_), .Y(_7333_) );
NOR2X1 NOR2X1_457 ( .A(_5358__bF_buf5), .B(_7333_), .Y(_7334_) );
INVX1 INVX1_589 ( .A(cpuregs_24_[28]), .Y(_7335_) );
NAND2X1 NAND2X1_443 ( .A(decoded_rs2_0_bF_buf69_), .B(cpuregs_25_[28]), .Y(_7336_) );
OAI21X1 OAI21X1_1127 ( .A(_7335_), .B(decoded_rs2_0_bF_buf68_), .C(_7336_), .Y(_7337_) );
INVX1 INVX1_590 ( .A(cpuregs_27_[28]), .Y(_7338_) );
OAI21X1 OAI21X1_1128 ( .A(decoded_rs2_0_bF_buf67_), .B(cpuregs_26_[28]), .C(decoded_rs2_1_bF_buf37_), .Y(_7339_) );
AOI21X1 AOI21X1_284 ( .A(decoded_rs2_0_bF_buf66_), .B(_7338_), .C(_7339_), .Y(_7340_) );
AOI21X1 AOI21X1_285 ( .A(_5349__bF_buf9), .B(_7337_), .C(_7340_), .Y(_7341_) );
NOR2X1 NOR2X1_458 ( .A(decoded_rs2_2_bF_buf2_), .B(_7341_), .Y(_7342_) );
OAI21X1 OAI21X1_1129 ( .A(_7334_), .B(_7342_), .C(decoded_rs2_4_bF_buf5_), .Y(_7343_) );
NOR2X1 NOR2X1_459 ( .A(cpuregs_8_[28]), .B(decoded_rs2_0_bF_buf65_), .Y(_7344_) );
OAI21X1 OAI21X1_1130 ( .A(_5362__bF_buf8), .B(cpuregs_9_[28]), .C(_5349__bF_buf8), .Y(_7345_) );
NOR2X1 NOR2X1_460 ( .A(cpuregs_11_[28]), .B(_5362__bF_buf7), .Y(_7346_) );
OAI21X1 OAI21X1_1131 ( .A(decoded_rs2_0_bF_buf64_), .B(cpuregs_10_[28]), .C(decoded_rs2_1_bF_buf36_), .Y(_7347_) );
OAI22X1 OAI22X1_78 ( .A(_7346_), .B(_7347_), .C(_7345_), .D(_7344_), .Y(_7348_) );
INVX1 INVX1_591 ( .A(cpuregs_13_[28]), .Y(_7349_) );
AOI21X1 AOI21X1_286 ( .A(decoded_rs2_0_bF_buf63_), .B(_7349_), .C(decoded_rs2_1_bF_buf35_), .Y(_7350_) );
OAI21X1 OAI21X1_1132 ( .A(decoded_rs2_0_bF_buf62_), .B(cpuregs_12_[28]), .C(_7350_), .Y(_7351_) );
NOR2X1 NOR2X1_461 ( .A(cpuregs_15_[28]), .B(_5362__bF_buf6), .Y(_7352_) );
OAI21X1 OAI21X1_1133 ( .A(decoded_rs2_0_bF_buf61_), .B(cpuregs_14_[28]), .C(decoded_rs2_1_bF_buf34_), .Y(_7353_) );
OAI21X1 OAI21X1_1134 ( .A(_7352_), .B(_7353_), .C(_7351_), .Y(_7354_) );
MUX2X1 MUX2X1_131 ( .A(_7354_), .B(_7348_), .S(decoded_rs2_2_bF_buf1_), .Y(_7355_) );
OAI21X1 OAI21X1_1135 ( .A(decoded_rs2_4_bF_buf4_), .B(_7355_), .C(_7343_), .Y(_7356_) );
AND2X2 AND2X2_45 ( .A(_7356_), .B(decoded_rs2_3_bF_buf1_), .Y(_7357_) );
OAI21X1 OAI21X1_1136 ( .A(_7357_), .B(_7326_), .C(_6422_), .Y(_7358_) );
AOI21X1 AOI21X1_287 ( .A(decoded_imm_28_), .B(_5849__bF_buf1), .C(_4540__bF_buf6), .Y(_7359_) );
AOI22X1 AOI22X1_41 ( .A(_5005_), .B(_4540__bF_buf5), .C(_7358_), .D(_7359_), .Y(_82__28_) );
NOR2X1 NOR2X1_462 ( .A(decoded_rs2_0_bF_buf60_), .B(cpuregs_0_[29]), .Y(_7360_) );
OAI21X1 OAI21X1_1137 ( .A(_5362__bF_buf5), .B(cpuregs_1_[29]), .C(_5349__bF_buf7), .Y(_7361_) );
NOR2X1 NOR2X1_463 ( .A(cpuregs_3_[29]), .B(_5362__bF_buf4), .Y(_7362_) );
OAI21X1 OAI21X1_1138 ( .A(decoded_rs2_0_bF_buf59_), .B(cpuregs_2_[29]), .C(decoded_rs2_1_bF_buf33_), .Y(_7363_) );
OAI22X1 OAI22X1_79 ( .A(_7362_), .B(_7363_), .C(_7361_), .D(_7360_), .Y(_7364_) );
NOR2X1 NOR2X1_464 ( .A(decoded_rs2_2_bF_buf0_), .B(_7364_), .Y(_7365_) );
NOR2X1 NOR2X1_465 ( .A(decoded_rs2_0_bF_buf58_), .B(cpuregs_4_[29]), .Y(_7366_) );
OAI21X1 OAI21X1_1139 ( .A(_5362__bF_buf3), .B(cpuregs_5_[29]), .C(_5349__bF_buf6), .Y(_7367_) );
NOR2X1 NOR2X1_466 ( .A(cpuregs_7_[29]), .B(_5362__bF_buf2), .Y(_7368_) );
OAI21X1 OAI21X1_1140 ( .A(cpuregs_6_[29]), .B(decoded_rs2_0_bF_buf57_), .C(decoded_rs2_1_bF_buf32_), .Y(_7369_) );
OAI22X1 OAI22X1_80 ( .A(_7368_), .B(_7369_), .C(_7367_), .D(_7366_), .Y(_7370_) );
OAI21X1 OAI21X1_1141 ( .A(_7370_), .B(_5358__bF_buf4), .C(_5348__bF_buf3), .Y(_7371_) );
INVX1 INVX1_592 ( .A(cpuregs_13_[29]), .Y(_7372_) );
AOI21X1 AOI21X1_288 ( .A(decoded_rs2_0_bF_buf56_), .B(_7372_), .C(decoded_rs2_1_bF_buf31_), .Y(_7373_) );
OAI21X1 OAI21X1_1142 ( .A(decoded_rs2_0_bF_buf55_), .B(cpuregs_12_[29]), .C(_7373_), .Y(_7374_) );
NOR2X1 NOR2X1_467 ( .A(cpuregs_15_[29]), .B(_5362__bF_buf1), .Y(_7375_) );
OAI21X1 OAI21X1_1143 ( .A(decoded_rs2_0_bF_buf54_), .B(cpuregs_14_[29]), .C(decoded_rs2_1_bF_buf30_), .Y(_7376_) );
OAI21X1 OAI21X1_1144 ( .A(_7375_), .B(_7376_), .C(_7374_), .Y(_7377_) );
NOR2X1 NOR2X1_468 ( .A(_5358__bF_buf3), .B(_7377_), .Y(_7378_) );
INVX1 INVX1_593 ( .A(cpuregs_9_[29]), .Y(_7379_) );
AOI21X1 AOI21X1_289 ( .A(decoded_rs2_0_bF_buf53_), .B(_7379_), .C(decoded_rs2_1_bF_buf29_), .Y(_7380_) );
OAI21X1 OAI21X1_1145 ( .A(cpuregs_8_[29]), .B(decoded_rs2_0_bF_buf52_), .C(_7380_), .Y(_7381_) );
NOR2X1 NOR2X1_469 ( .A(cpuregs_11_[29]), .B(_5362__bF_buf0), .Y(_7382_) );
OAI21X1 OAI21X1_1146 ( .A(decoded_rs2_0_bF_buf51_), .B(cpuregs_10_[29]), .C(decoded_rs2_1_bF_buf28_), .Y(_7383_) );
OAI21X1 OAI21X1_1147 ( .A(_7382_), .B(_7383_), .C(_7381_), .Y(_7384_) );
OAI21X1 OAI21X1_1148 ( .A(_7384_), .B(decoded_rs2_2_bF_buf8_), .C(decoded_rs2_3_bF_buf0_), .Y(_7385_) );
OAI22X1 OAI22X1_81 ( .A(_7365_), .B(_7371_), .C(_7385_), .D(_7378_), .Y(_7386_) );
INVX1 INVX1_594 ( .A(cpuregs_26_[29]), .Y(_7387_) );
OAI21X1 OAI21X1_1149 ( .A(_7387_), .B(decoded_rs2_0_bF_buf50_), .C(decoded_rs2_1_bF_buf27_), .Y(_7388_) );
AOI21X1 AOI21X1_290 ( .A(decoded_rs2_0_bF_buf49_), .B(cpuregs_27_[29]), .C(_7388_), .Y(_7389_) );
AND2X2 AND2X2_46 ( .A(decoded_rs2_0_bF_buf48_), .B(cpuregs_25_[29]), .Y(_7390_) );
INVX1 INVX1_595 ( .A(cpuregs_24_[29]), .Y(_7391_) );
OAI21X1 OAI21X1_1150 ( .A(_7391_), .B(decoded_rs2_0_bF_buf47_), .C(_5349__bF_buf5), .Y(_7392_) );
OAI21X1 OAI21X1_1151 ( .A(_7392_), .B(_7390_), .C(_5358__bF_buf2), .Y(_7393_) );
INVX1 INVX1_596 ( .A(cpuregs_28_[29]), .Y(_7394_) );
NAND2X1 NAND2X1_444 ( .A(decoded_rs2_0_bF_buf46_), .B(cpuregs_29_[29]), .Y(_7395_) );
OAI21X1 OAI21X1_1152 ( .A(_7394_), .B(decoded_rs2_0_bF_buf45_), .C(_7395_), .Y(_7396_) );
INVX1 INVX1_597 ( .A(cpuregs_30_[29]), .Y(_7397_) );
NAND2X1 NAND2X1_445 ( .A(decoded_rs2_0_bF_buf44_), .B(cpuregs_31_[29]), .Y(_7398_) );
OAI21X1 OAI21X1_1153 ( .A(_7397_), .B(decoded_rs2_0_bF_buf43_), .C(_7398_), .Y(_7399_) );
MUX2X1 MUX2X1_132 ( .A(_7399_), .B(_7396_), .S(decoded_rs2_1_bF_buf26_), .Y(_7400_) );
OAI22X1 OAI22X1_82 ( .A(_7393_), .B(_7389_), .C(_7400_), .D(_5358__bF_buf1), .Y(_7401_) );
INVX1 INVX1_598 ( .A(cpuregs_16_[29]), .Y(_7402_) );
NAND2X1 NAND2X1_446 ( .A(decoded_rs2_0_bF_buf42_), .B(cpuregs_17_[29]), .Y(_7403_) );
OAI21X1 OAI21X1_1154 ( .A(_7402_), .B(decoded_rs2_0_bF_buf41_), .C(_7403_), .Y(_7404_) );
INVX1 INVX1_599 ( .A(cpuregs_19_[29]), .Y(_7405_) );
OAI21X1 OAI21X1_1155 ( .A(decoded_rs2_0_bF_buf40_), .B(cpuregs_18_[29]), .C(decoded_rs2_1_bF_buf25_), .Y(_7406_) );
AOI21X1 AOI21X1_291 ( .A(decoded_rs2_0_bF_buf39_), .B(_7405_), .C(_7406_), .Y(_7407_) );
AOI21X1 AOI21X1_292 ( .A(_5349__bF_buf4), .B(_7404_), .C(_7407_), .Y(_7408_) );
NAND2X1 NAND2X1_447 ( .A(_5358__bF_buf0), .B(_7408_), .Y(_7409_) );
INVX1 INVX1_600 ( .A(cpuregs_20_[29]), .Y(_7410_) );
NAND2X1 NAND2X1_448 ( .A(decoded_rs2_0_bF_buf38_), .B(cpuregs_21_[29]), .Y(_7411_) );
OAI21X1 OAI21X1_1156 ( .A(_7410_), .B(decoded_rs2_0_bF_buf37_), .C(_7411_), .Y(_7412_) );
INVX1 INVX1_601 ( .A(cpuregs_22_[29]), .Y(_7413_) );
NAND2X1 NAND2X1_449 ( .A(decoded_rs2_0_bF_buf36_), .B(cpuregs_23_[29]), .Y(_7414_) );
OAI21X1 OAI21X1_1157 ( .A(_7413_), .B(decoded_rs2_0_bF_buf35_), .C(_7414_), .Y(_7415_) );
MUX2X1 MUX2X1_133 ( .A(_7415_), .B(_7412_), .S(decoded_rs2_1_bF_buf24_), .Y(_7416_) );
AOI21X1 AOI21X1_293 ( .A(decoded_rs2_2_bF_buf7_), .B(_7416_), .C(decoded_rs2_3_bF_buf6_), .Y(_7417_) );
AOI22X1 AOI22X1_42 ( .A(_7417_), .B(_7409_), .C(decoded_rs2_3_bF_buf5_), .D(_7401_), .Y(_7418_) );
AOI21X1 AOI21X1_294 ( .A(decoded_rs2_4_bF_buf3_), .B(_7418_), .C(_5890__bF_buf1), .Y(_7419_) );
OAI21X1 OAI21X1_1158 ( .A(decoded_rs2_4_bF_buf2_), .B(_7386_), .C(_7419_), .Y(_7420_) );
AOI21X1 AOI21X1_295 ( .A(decoded_imm_29_), .B(_5849__bF_buf0), .C(_4540__bF_buf4), .Y(_7421_) );
AOI22X1 AOI22X1_43 ( .A(_5010_), .B(_4540__bF_buf3), .C(_7420_), .D(_7421_), .Y(_82__29_) );
INVX1 INVX1_602 ( .A(cpuregs_20_[30]), .Y(_7422_) );
OAI21X1 OAI21X1_1159 ( .A(_5358__bF_buf12), .B(_7422_), .C(_5362__bF_buf14), .Y(_7423_) );
AOI21X1 AOI21X1_296 ( .A(_5358__bF_buf11), .B(cpuregs_16_[30]), .C(_7423_), .Y(_7424_) );
INVX1 INVX1_603 ( .A(cpuregs_21_[30]), .Y(_7425_) );
OAI21X1 OAI21X1_1160 ( .A(_5358__bF_buf10), .B(_7425_), .C(decoded_rs2_0_bF_buf34_), .Y(_7426_) );
AOI21X1 AOI21X1_297 ( .A(_5358__bF_buf9), .B(cpuregs_17_[30]), .C(_7426_), .Y(_7427_) );
OAI21X1 OAI21X1_1161 ( .A(_7424_), .B(_7427_), .C(_5349__bF_buf3), .Y(_7428_) );
INVX1 INVX1_604 ( .A(cpuregs_22_[30]), .Y(_7429_) );
OAI21X1 OAI21X1_1162 ( .A(_5358__bF_buf8), .B(_7429_), .C(_5362__bF_buf13), .Y(_7430_) );
AOI21X1 AOI21X1_298 ( .A(_5358__bF_buf7), .B(cpuregs_18_[30]), .C(_7430_), .Y(_7431_) );
INVX1 INVX1_605 ( .A(cpuregs_23_[30]), .Y(_7432_) );
OAI21X1 OAI21X1_1163 ( .A(_5358__bF_buf6), .B(_7432_), .C(decoded_rs2_0_bF_buf33_), .Y(_7433_) );
AOI21X1 AOI21X1_299 ( .A(_5358__bF_buf5), .B(cpuregs_19_[30]), .C(_7433_), .Y(_7434_) );
OAI21X1 OAI21X1_1164 ( .A(_7431_), .B(_7434_), .C(decoded_rs2_1_bF_buf23_), .Y(_7435_) );
NAND3X1 NAND3X1_31 ( .A(decoded_rs2_4_bF_buf1_), .B(_7428_), .C(_7435_), .Y(_7436_) );
INVX1 INVX1_606 ( .A(cpuregs_6_[30]), .Y(_7437_) );
AOI21X1 AOI21X1_300 ( .A(decoded_rs2_1_bF_buf22_), .B(_7437_), .C(decoded_rs2_0_bF_buf32_), .Y(_7438_) );
OAI21X1 OAI21X1_1165 ( .A(decoded_rs2_1_bF_buf21_), .B(cpuregs_4_[30]), .C(_7438_), .Y(_7439_) );
NOR2X1 NOR2X1_470 ( .A(cpuregs_5_[30]), .B(decoded_rs2_1_bF_buf20_), .Y(_7440_) );
OAI21X1 OAI21X1_1166 ( .A(_5349__bF_buf2), .B(cpuregs_7_[30]), .C(decoded_rs2_0_bF_buf31_), .Y(_7441_) );
OAI21X1 OAI21X1_1167 ( .A(_7440_), .B(_7441_), .C(_7439_), .Y(_7442_) );
INVX1 INVX1_607 ( .A(cpuregs_2_[30]), .Y(_7443_) );
AOI21X1 AOI21X1_301 ( .A(decoded_rs2_1_bF_buf19_), .B(_7443_), .C(decoded_rs2_0_bF_buf30_), .Y(_7444_) );
OAI21X1 OAI21X1_1168 ( .A(decoded_rs2_1_bF_buf18_), .B(cpuregs_0_[30]), .C(_7444_), .Y(_7445_) );
NOR2X1 NOR2X1_471 ( .A(decoded_rs2_1_bF_buf17_), .B(cpuregs_1_[30]), .Y(_7446_) );
OAI21X1 OAI21X1_1169 ( .A(_5349__bF_buf1), .B(cpuregs_3_[30]), .C(decoded_rs2_0_bF_buf29_), .Y(_7447_) );
OAI21X1 OAI21X1_1170 ( .A(_7446_), .B(_7447_), .C(_7445_), .Y(_7448_) );
MUX2X1 MUX2X1_134 ( .A(_7448_), .B(_7442_), .S(_5358__bF_buf4), .Y(_7449_) );
OAI21X1 OAI21X1_1171 ( .A(decoded_rs2_4_bF_buf0_), .B(_7449_), .C(_7436_), .Y(_7450_) );
AND2X2 AND2X2_47 ( .A(_7450_), .B(_5348__bF_buf2), .Y(_7451_) );
INVX1 INVX1_608 ( .A(cpuregs_29_[30]), .Y(_7452_) );
NAND2X1 NAND2X1_450 ( .A(decoded_rs2_1_bF_buf16_), .B(cpuregs_31_[30]), .Y(_7453_) );
OAI21X1 OAI21X1_1172 ( .A(_7452_), .B(decoded_rs2_1_bF_buf15_), .C(_7453_), .Y(_7454_) );
INVX1 INVX1_609 ( .A(cpuregs_28_[30]), .Y(_7455_) );
NAND2X1 NAND2X1_451 ( .A(decoded_rs2_1_bF_buf14_), .B(cpuregs_30_[30]), .Y(_7456_) );
OAI21X1 OAI21X1_1173 ( .A(_7455_), .B(decoded_rs2_1_bF_buf13_), .C(_7456_), .Y(_7457_) );
MUX2X1 MUX2X1_135 ( .A(_7457_), .B(_7454_), .S(_5362__bF_buf12), .Y(_7458_) );
NOR2X1 NOR2X1_472 ( .A(_5358__bF_buf3), .B(_7458_), .Y(_7459_) );
INVX1 INVX1_610 ( .A(cpuregs_24_[30]), .Y(_7460_) );
NAND2X1 NAND2X1_452 ( .A(decoded_rs2_0_bF_buf28_), .B(cpuregs_25_[30]), .Y(_7461_) );
OAI21X1 OAI21X1_1174 ( .A(_7460_), .B(decoded_rs2_0_bF_buf27_), .C(_7461_), .Y(_7462_) );
INVX1 INVX1_611 ( .A(cpuregs_27_[30]), .Y(_7463_) );
OAI21X1 OAI21X1_1175 ( .A(decoded_rs2_0_bF_buf26_), .B(cpuregs_26_[30]), .C(decoded_rs2_1_bF_buf12_), .Y(_7464_) );
AOI21X1 AOI21X1_302 ( .A(decoded_rs2_0_bF_buf25_), .B(_7463_), .C(_7464_), .Y(_7465_) );
AOI21X1 AOI21X1_303 ( .A(_5349__bF_buf0), .B(_7462_), .C(_7465_), .Y(_7466_) );
NOR2X1 NOR2X1_473 ( .A(decoded_rs2_2_bF_buf6_), .B(_7466_), .Y(_7467_) );
OAI21X1 OAI21X1_1176 ( .A(_7459_), .B(_7467_), .C(decoded_rs2_4_bF_buf7_), .Y(_7468_) );
NOR2X1 NOR2X1_474 ( .A(cpuregs_8_[30]), .B(decoded_rs2_0_bF_buf24_), .Y(_7469_) );
OAI21X1 OAI21X1_1177 ( .A(_5362__bF_buf11), .B(cpuregs_9_[30]), .C(_5349__bF_buf11), .Y(_7470_) );
NOR2X1 NOR2X1_475 ( .A(cpuregs_11_[30]), .B(_5362__bF_buf10), .Y(_7471_) );
OAI21X1 OAI21X1_1178 ( .A(decoded_rs2_0_bF_buf23_), .B(cpuregs_10_[30]), .C(decoded_rs2_1_bF_buf11_), .Y(_7472_) );
OAI22X1 OAI22X1_83 ( .A(_7471_), .B(_7472_), .C(_7470_), .D(_7469_), .Y(_7473_) );
NOR2X1 NOR2X1_476 ( .A(decoded_rs2_0_bF_buf22_), .B(cpuregs_12_[30]), .Y(_7474_) );
OAI21X1 OAI21X1_1179 ( .A(_5362__bF_buf9), .B(cpuregs_13_[30]), .C(_5349__bF_buf10), .Y(_7475_) );
NOR2X1 NOR2X1_477 ( .A(cpuregs_15_[30]), .B(_5362__bF_buf8), .Y(_7476_) );
OAI21X1 OAI21X1_1180 ( .A(decoded_rs2_0_bF_buf21_), .B(cpuregs_14_[30]), .C(decoded_rs2_1_bF_buf10_), .Y(_7477_) );
OAI22X1 OAI22X1_84 ( .A(_7476_), .B(_7477_), .C(_7475_), .D(_7474_), .Y(_7478_) );
MUX2X1 MUX2X1_136 ( .A(_7478_), .B(_7473_), .S(decoded_rs2_2_bF_buf5_), .Y(_7479_) );
OAI21X1 OAI21X1_1181 ( .A(decoded_rs2_4_bF_buf6_), .B(_7479_), .C(_7468_), .Y(_7480_) );
AND2X2 AND2X2_48 ( .A(_7480_), .B(decoded_rs2_3_bF_buf4_), .Y(_7481_) );
OAI21X1 OAI21X1_1182 ( .A(_7481_), .B(_7451_), .C(_6422_), .Y(_7482_) );
AOI21X1 AOI21X1_304 ( .A(decoded_imm_30_), .B(_5849__bF_buf4), .C(_4540__bF_buf2), .Y(_7483_) );
AOI22X1 AOI22X1_44 ( .A(_4999_), .B(_4540__bF_buf1), .C(_7482_), .D(_7483_), .Y(_82__30_) );
INVX1 INVX1_612 ( .A(cpuregs_0_[31]), .Y(_7484_) );
NAND2X1 NAND2X1_453 ( .A(decoded_rs2_0_bF_buf20_), .B(cpuregs_1_[31]), .Y(_7485_) );
OAI21X1 OAI21X1_1183 ( .A(_7484_), .B(decoded_rs2_0_bF_buf19_), .C(_7485_), .Y(_7486_) );
INVX1 INVX1_613 ( .A(cpuregs_2_[31]), .Y(_7487_) );
NAND2X1 NAND2X1_454 ( .A(decoded_rs2_0_bF_buf18_), .B(cpuregs_3_[31]), .Y(_7488_) );
OAI21X1 OAI21X1_1184 ( .A(_7487_), .B(decoded_rs2_0_bF_buf17_), .C(_7488_), .Y(_7489_) );
MUX2X1 MUX2X1_137 ( .A(_7489_), .B(_7486_), .S(decoded_rs2_1_bF_buf9_), .Y(_7490_) );
NAND2X1 NAND2X1_455 ( .A(_5358__bF_buf2), .B(_7490_), .Y(_7491_) );
NOR2X1 NOR2X1_478 ( .A(decoded_rs2_0_bF_buf16_), .B(cpuregs_4_[31]), .Y(_7492_) );
OAI21X1 OAI21X1_1185 ( .A(_5362__bF_buf7), .B(cpuregs_5_[31]), .C(_5349__bF_buf9), .Y(_7493_) );
NOR2X1 NOR2X1_479 ( .A(cpuregs_7_[31]), .B(_5362__bF_buf6), .Y(_7494_) );
OAI21X1 OAI21X1_1186 ( .A(cpuregs_6_[31]), .B(decoded_rs2_0_bF_buf15_), .C(decoded_rs2_1_bF_buf8_), .Y(_7495_) );
OAI22X1 OAI22X1_85 ( .A(_7494_), .B(_7495_), .C(_7493_), .D(_7492_), .Y(_7496_) );
OAI21X1 OAI21X1_1187 ( .A(_5358__bF_buf1), .B(_7496_), .C(_7491_), .Y(_7497_) );
INVX1 INVX1_614 ( .A(cpuregs_9_[31]), .Y(_7498_) );
NAND2X1 NAND2X1_456 ( .A(cpuregs_8_[31]), .B(_5362__bF_buf5), .Y(_7499_) );
OAI21X1 OAI21X1_1188 ( .A(_5362__bF_buf4), .B(_7498_), .C(_7499_), .Y(_7500_) );
INVX1 INVX1_615 ( .A(cpuregs_11_[31]), .Y(_7501_) );
NAND2X1 NAND2X1_457 ( .A(cpuregs_10_[31]), .B(_5362__bF_buf3), .Y(_7502_) );
OAI21X1 OAI21X1_1189 ( .A(_5362__bF_buf2), .B(_7501_), .C(_7502_), .Y(_7503_) );
MUX2X1 MUX2X1_138 ( .A(_7503_), .B(_7500_), .S(decoded_rs2_1_bF_buf7_), .Y(_7504_) );
INVX1 INVX1_616 ( .A(cpuregs_13_[31]), .Y(_7505_) );
OAI21X1 OAI21X1_1190 ( .A(_7505_), .B(decoded_rs2_1_bF_buf6_), .C(decoded_rs2_0_bF_buf14_), .Y(_7506_) );
AOI21X1 AOI21X1_305 ( .A(decoded_rs2_1_bF_buf5_), .B(cpuregs_15_[31]), .C(_7506_), .Y(_7507_) );
INVX1 INVX1_617 ( .A(cpuregs_14_[31]), .Y(_7508_) );
NOR2X1 NOR2X1_480 ( .A(_5349__bF_buf8), .B(_7508_), .Y(_7509_) );
INVX1 INVX1_618 ( .A(cpuregs_12_[31]), .Y(_7510_) );
OAI21X1 OAI21X1_1191 ( .A(_7510_), .B(decoded_rs2_1_bF_buf4_), .C(_5362__bF_buf1), .Y(_7511_) );
OAI21X1 OAI21X1_1192 ( .A(_7511_), .B(_7509_), .C(decoded_rs2_2_bF_buf4_), .Y(_7512_) );
OAI22X1 OAI22X1_86 ( .A(_7512_), .B(_7507_), .C(_7504_), .D(decoded_rs2_2_bF_buf3_), .Y(_7513_) );
NAND2X1 NAND2X1_458 ( .A(decoded_rs2_3_bF_buf3_), .B(_7513_), .Y(_7514_) );
OAI21X1 OAI21X1_1193 ( .A(_7497_), .B(decoded_rs2_3_bF_buf2_), .C(_7514_), .Y(_7515_) );
INVX1 INVX1_619 ( .A(cpuregs_16_[31]), .Y(_7516_) );
NAND2X1 NAND2X1_459 ( .A(decoded_rs2_0_bF_buf13_), .B(cpuregs_17_[31]), .Y(_7517_) );
OAI21X1 OAI21X1_1194 ( .A(_7516_), .B(decoded_rs2_0_bF_buf12_), .C(_7517_), .Y(_7518_) );
INVX1 INVX1_620 ( .A(cpuregs_18_[31]), .Y(_7519_) );
NAND2X1 NAND2X1_460 ( .A(decoded_rs2_0_bF_buf11_), .B(cpuregs_19_[31]), .Y(_7520_) );
OAI21X1 OAI21X1_1195 ( .A(_7519_), .B(decoded_rs2_0_bF_buf10_), .C(_7520_), .Y(_7521_) );
MUX2X1 MUX2X1_139 ( .A(_7521_), .B(_7518_), .S(decoded_rs2_1_bF_buf3_), .Y(_7522_) );
INVX1 INVX1_621 ( .A(cpuregs_20_[31]), .Y(_7523_) );
NAND2X1 NAND2X1_461 ( .A(decoded_rs2_0_bF_buf9_), .B(cpuregs_21_[31]), .Y(_7524_) );
OAI21X1 OAI21X1_1196 ( .A(_7523_), .B(decoded_rs2_0_bF_buf8_), .C(_7524_), .Y(_7525_) );
INVX1 INVX1_622 ( .A(cpuregs_22_[31]), .Y(_7526_) );
NAND2X1 NAND2X1_462 ( .A(decoded_rs2_0_bF_buf7_), .B(cpuregs_23_[31]), .Y(_7527_) );
OAI21X1 OAI21X1_1197 ( .A(_7526_), .B(decoded_rs2_0_bF_buf6_), .C(_7527_), .Y(_7528_) );
MUX2X1 MUX2X1_140 ( .A(_7528_), .B(_7525_), .S(decoded_rs2_1_bF_buf2_), .Y(_7529_) );
MUX2X1 MUX2X1_141 ( .A(_7529_), .B(_7522_), .S(decoded_rs2_2_bF_buf2_), .Y(_7530_) );
INVX1 INVX1_623 ( .A(cpuregs_26_[31]), .Y(_7531_) );
OAI21X1 OAI21X1_1198 ( .A(_7531_), .B(decoded_rs2_0_bF_buf5_), .C(decoded_rs2_1_bF_buf1_), .Y(_7532_) );
AOI21X1 AOI21X1_306 ( .A(decoded_rs2_0_bF_buf4_), .B(cpuregs_27_[31]), .C(_7532_), .Y(_7533_) );
AND2X2 AND2X2_49 ( .A(decoded_rs2_0_bF_buf3_), .B(cpuregs_25_[31]), .Y(_7534_) );
INVX1 INVX1_624 ( .A(cpuregs_24_[31]), .Y(_7535_) );
OAI21X1 OAI21X1_1199 ( .A(_7535_), .B(decoded_rs2_0_bF_buf2_), .C(_5349__bF_buf7), .Y(_7536_) );
OAI21X1 OAI21X1_1200 ( .A(_7536_), .B(_7534_), .C(_5358__bF_buf0), .Y(_7537_) );
INVX1 INVX1_625 ( .A(cpuregs_28_[31]), .Y(_7538_) );
NAND2X1 NAND2X1_463 ( .A(decoded_rs2_0_bF_buf1_), .B(cpuregs_29_[31]), .Y(_7539_) );
OAI21X1 OAI21X1_1201 ( .A(_7538_), .B(decoded_rs2_0_bF_buf0_), .C(_7539_), .Y(_7540_) );
INVX1 INVX1_626 ( .A(cpuregs_30_[31]), .Y(_7541_) );
NAND2X1 NAND2X1_464 ( .A(decoded_rs2_0_bF_buf78_), .B(cpuregs_31_[31]), .Y(_7542_) );
OAI21X1 OAI21X1_1202 ( .A(_7541_), .B(decoded_rs2_0_bF_buf77_), .C(_7542_), .Y(_7543_) );
MUX2X1 MUX2X1_142 ( .A(_7543_), .B(_7540_), .S(decoded_rs2_1_bF_buf0_), .Y(_7544_) );
OAI22X1 OAI22X1_87 ( .A(_7537_), .B(_7533_), .C(_7544_), .D(_5358__bF_buf12), .Y(_7545_) );
MUX2X1 MUX2X1_143 ( .A(_7545_), .B(_7530_), .S(decoded_rs2_3_bF_buf1_), .Y(_7546_) );
AOI21X1 AOI21X1_307 ( .A(decoded_rs2_4_bF_buf5_), .B(_7546_), .C(_5890__bF_buf0), .Y(_7547_) );
OAI21X1 OAI21X1_1203 ( .A(_7515_), .B(decoded_rs2_4_bF_buf4_), .C(_7547_), .Y(_7548_) );
AOI21X1 AOI21X1_308 ( .A(decoded_imm_31_), .B(_5849__bF_buf3), .C(_4540__bF_buf0), .Y(_7549_) );
AOI22X1 AOI22X1_45 ( .A(_4994_), .B(_4540__bF_buf6), .C(_7548_), .D(_7549_), .Y(_82__31_) );
INVX1 INVX1_627 ( .A(is_lui_auipc_jal), .Y(_7550_) );
NOR2X1 NOR2X1_481 ( .A(instr_lui), .B(_7550_), .Y(_7551_) );
INVX1 INVX1_628 ( .A(decoded_rs1_4_bF_buf4_), .Y(_7552_) );
AOI21X1 AOI21X1_309 ( .A(decoded_rs1_1_bF_buf44_), .B(_5404_), .C(decoded_rs1_0_bF_buf57_), .Y(_7553_) );
OAI21X1 OAI21X1_1204 ( .A(cpuregs_16_[0]), .B(decoded_rs1_1_bF_buf43_), .C(_7553_), .Y(_7554_) );
NOR2X1 NOR2X1_482 ( .A(cpuregs_17_[0]), .B(decoded_rs1_1_bF_buf42_), .Y(_7555_) );
INVX1 INVX1_629 ( .A(decoded_rs1_1_bF_buf41_), .Y(_7556_) );
OAI21X1 OAI21X1_1205 ( .A(_7556__bF_buf42), .B(cpuregs_19_[0]), .C(decoded_rs1_0_bF_buf56_), .Y(_7557_) );
OAI21X1 OAI21X1_1206 ( .A(_7555_), .B(_7557_), .C(_7554_), .Y(_7558_) );
NOR2X1 NOR2X1_483 ( .A(decoded_rs1_2_bF_buf12_), .B(_7558_), .Y(_7559_) );
INVX1 INVX1_630 ( .A(decoded_rs1_2_bF_buf11_), .Y(_7560_) );
INVX1 INVX1_631 ( .A(decoded_rs1_3_bF_buf6_), .Y(_7561_) );
AOI21X1 AOI21X1_310 ( .A(decoded_rs1_1_bF_buf40_), .B(_5411_), .C(decoded_rs1_0_bF_buf55_), .Y(_7562_) );
OAI21X1 OAI21X1_1207 ( .A(cpuregs_20_[0]), .B(decoded_rs1_1_bF_buf39_), .C(_7562_), .Y(_7563_) );
NOR2X1 NOR2X1_484 ( .A(cpuregs_21_[0]), .B(decoded_rs1_1_bF_buf38_), .Y(_7564_) );
OAI21X1 OAI21X1_1208 ( .A(_7556__bF_buf41), .B(cpuregs_23_[0]), .C(decoded_rs1_0_bF_buf54_), .Y(_7565_) );
OAI21X1 OAI21X1_1209 ( .A(_7564_), .B(_7565_), .C(_7563_), .Y(_7566_) );
OAI21X1 OAI21X1_1210 ( .A(_7566_), .B(_7560__bF_buf12), .C(_7561__bF_buf6), .Y(_7567_) );
NOR2X1 NOR2X1_485 ( .A(cpuregs_24_[0]), .B(decoded_rs1_0_bF_buf53_), .Y(_7568_) );
INVX1 INVX1_632 ( .A(decoded_rs1_0_bF_buf52_), .Y(_7569_) );
OAI21X1 OAI21X1_1211 ( .A(_7569__bF_buf48), .B(cpuregs_25_[0]), .C(_7556__bF_buf40), .Y(_7570_) );
NOR2X1 NOR2X1_486 ( .A(cpuregs_27_[0]), .B(_7569__bF_buf47), .Y(_7571_) );
OAI21X1 OAI21X1_1212 ( .A(cpuregs_26_[0]), .B(decoded_rs1_0_bF_buf51_), .C(decoded_rs1_1_bF_buf37_), .Y(_7572_) );
OAI22X1 OAI22X1_88 ( .A(_7571_), .B(_7572_), .C(_7570_), .D(_7568_), .Y(_7573_) );
NOR2X1 NOR2X1_487 ( .A(decoded_rs1_2_bF_buf10_), .B(_7573_), .Y(_7574_) );
NOR2X1 NOR2X1_488 ( .A(cpuregs_28_[0]), .B(decoded_rs1_0_bF_buf50_), .Y(_7575_) );
OAI21X1 OAI21X1_1213 ( .A(_7569__bF_buf46), .B(cpuregs_29_[0]), .C(_7556__bF_buf39), .Y(_7576_) );
NOR2X1 NOR2X1_489 ( .A(cpuregs_31_[0]), .B(_7569__bF_buf45), .Y(_7577_) );
OAI21X1 OAI21X1_1214 ( .A(cpuregs_30_[0]), .B(decoded_rs1_0_bF_buf49_), .C(decoded_rs1_1_bF_buf36_), .Y(_7578_) );
OAI22X1 OAI22X1_89 ( .A(_7577_), .B(_7578_), .C(_7576_), .D(_7575_), .Y(_7579_) );
OAI21X1 OAI21X1_1215 ( .A(_7579_), .B(_7560__bF_buf11), .C(decoded_rs1_3_bF_buf5_), .Y(_7580_) );
OAI22X1 OAI22X1_90 ( .A(_7574_), .B(_7580_), .C(_7567_), .D(_7559_), .Y(_7581_) );
NOR2X1 NOR2X1_490 ( .A(_7552__bF_buf5), .B(_7581_), .Y(_7582_) );
NOR2X1 NOR2X1_491 ( .A(decoded_rs1_4_bF_buf3_), .B(decoded_rs1_0_bF_buf48_), .Y(_7583_) );
INVX1 INVX1_633 ( .A(_7583_), .Y(_7584_) );
NAND3X1 NAND3X1_32 ( .A(_7556__bF_buf38), .B(_7560__bF_buf10), .C(_7561__bF_buf5), .Y(_7585_) );
OAI21X1 OAI21X1_1216 ( .A(_7585_), .B(_7584_), .C(_7550_), .Y(_7586_) );
INVX1 INVX1_634 ( .A(_7586__bF_buf3), .Y(_7587_) );
AOI21X1 AOI21X1_311 ( .A(cpuregs_10_[0]), .B(_7569__bF_buf44), .C(_7556__bF_buf37), .Y(_7588_) );
OAI21X1 OAI21X1_1217 ( .A(_5363_), .B(_7569__bF_buf43), .C(_7588_), .Y(_7589_) );
OAI21X1 OAI21X1_1218 ( .A(_5359_), .B(decoded_rs1_0_bF_buf47_), .C(_7556__bF_buf36), .Y(_7590_) );
AOI21X1 AOI21X1_312 ( .A(cpuregs_9_[0]), .B(decoded_rs1_0_bF_buf46_), .C(_7590_), .Y(_7591_) );
NOR2X1 NOR2X1_492 ( .A(decoded_rs1_2_bF_buf9_), .B(_7591_), .Y(_7592_) );
NOR2X1 NOR2X1_493 ( .A(cpuregs_12_[0]), .B(decoded_rs1_0_bF_buf45_), .Y(_7593_) );
OAI21X1 OAI21X1_1219 ( .A(_7569__bF_buf42), .B(cpuregs_13_[0]), .C(_7556__bF_buf35), .Y(_7594_) );
NOR2X1 NOR2X1_494 ( .A(cpuregs_15_[0]), .B(_7569__bF_buf41), .Y(_7595_) );
OAI21X1 OAI21X1_1220 ( .A(cpuregs_14_[0]), .B(decoded_rs1_0_bF_buf44_), .C(decoded_rs1_1_bF_buf35_), .Y(_7596_) );
OAI22X1 OAI22X1_91 ( .A(_7595_), .B(_7596_), .C(_7594_), .D(_7593_), .Y(_7597_) );
AOI22X1 AOI22X1_46 ( .A(decoded_rs1_2_bF_buf8_), .B(_7597_), .C(_7592_), .D(_7589_), .Y(_7598_) );
NOR2X1 NOR2X1_495 ( .A(cpuregs_0_[0]), .B(decoded_rs1_0_bF_buf43_), .Y(_7599_) );
OAI21X1 OAI21X1_1221 ( .A(_7569__bF_buf40), .B(cpuregs_1_[0]), .C(_7556__bF_buf34), .Y(_7600_) );
NOR2X1 NOR2X1_496 ( .A(cpuregs_3_[0]), .B(_7569__bF_buf39), .Y(_7601_) );
OAI21X1 OAI21X1_1222 ( .A(cpuregs_2_[0]), .B(decoded_rs1_0_bF_buf42_), .C(decoded_rs1_1_bF_buf34_), .Y(_7602_) );
OAI22X1 OAI22X1_92 ( .A(_7601_), .B(_7602_), .C(_7600_), .D(_7599_), .Y(_7603_) );
NOR2X1 NOR2X1_497 ( .A(decoded_rs1_2_bF_buf7_), .B(_7603_), .Y(_7604_) );
NOR2X1 NOR2X1_498 ( .A(cpuregs_4_[0]), .B(decoded_rs1_0_bF_buf41_), .Y(_7605_) );
OAI21X1 OAI21X1_1223 ( .A(_7569__bF_buf38), .B(cpuregs_5_[0]), .C(_7556__bF_buf33), .Y(_7606_) );
NOR2X1 NOR2X1_499 ( .A(cpuregs_7_[0]), .B(_7569__bF_buf37), .Y(_7607_) );
OAI21X1 OAI21X1_1224 ( .A(cpuregs_6_[0]), .B(decoded_rs1_0_bF_buf40_), .C(decoded_rs1_1_bF_buf33_), .Y(_7608_) );
OAI22X1 OAI22X1_93 ( .A(_7607_), .B(_7608_), .C(_7606_), .D(_7605_), .Y(_7609_) );
OAI21X1 OAI21X1_1225 ( .A(_7609_), .B(_7560__bF_buf9), .C(_7561__bF_buf4), .Y(_7610_) );
OAI22X1 OAI22X1_94 ( .A(_7610_), .B(_7604_), .C(_7598_), .D(_7561__bF_buf3), .Y(_7611_) );
OAI21X1 OAI21X1_1226 ( .A(_7611_), .B(decoded_rs1_4_bF_buf2_), .C(_7587_), .Y(_7612_) );
NOR2X1 NOR2X1_500 ( .A(_7582_), .B(_7612_), .Y(_7613_) );
AOI21X1 AOI21X1_313 ( .A(reg_pc_0_), .B(_7551__bF_buf3), .C(_7613_), .Y(_7614_) );
NOR2X1 NOR2X1_501 ( .A(instr_srli), .B(instr_srl), .Y(_7615_) );
OAI21X1 OAI21X1_1227 ( .A(instr_slli), .B(instr_sll), .C(_7615_), .Y(_7616_) );
OAI21X1 OAI21X1_1228 ( .A(_4580__bF_buf2), .B(_10734__1_), .C(_7616_), .Y(_7617_) );
AOI21X1 AOI21X1_314 ( .A(_5180_), .B(_4580__bF_buf1), .C(_7617_), .Y(_7618_) );
NOR2X1 NOR2X1_502 ( .A(_10734__0_), .B(decoded_imm_0_), .Y(_7619_) );
INVX1 INVX1_635 ( .A(decoded_imm_0_), .Y(_7620_) );
NOR2X1 NOR2X1_503 ( .A(_4491_), .B(_7620_), .Y(_7621_) );
NOR2X1 NOR2X1_504 ( .A(_7619_), .B(_7621_), .Y(_7622_) );
OAI21X1 OAI21X1_1229 ( .A(_4442_), .B(_4430_), .C(_4435_), .Y(_7623_) );
INVX1 INVX1_636 ( .A(_7623__bF_buf4), .Y(_7624_) );
NOR2X1 NOR2X1_505 ( .A(cpu_state_3_bF_buf3_), .B(cpu_state_1_bF_buf1_), .Y(_7625_) );
INVX1 INVX1_637 ( .A(_7625_), .Y(_7626_) );
NOR2X1 NOR2X1_506 ( .A(cpu_state_0_), .B(_7626_), .Y(_7627_) );
NOR2X1 NOR2X1_507 ( .A(cpu_state_5_bF_buf1_), .B(_4446_), .Y(_7628_) );
NAND2X1 NAND2X1_465 ( .A(_7627_), .B(_7628_), .Y(_7629_) );
INVX1 INVX1_638 ( .A(_7629__bF_buf3), .Y(_7630_) );
OAI21X1 OAI21X1_1230 ( .A(_4442_), .B(_4430_), .C(_4427_), .Y(_7631_) );
INVX1 INVX1_639 ( .A(_7631__bF_buf5), .Y(_7632_) );
AOI22X1 AOI22X1_47 ( .A(_7624__bF_buf4), .B(cpu_state_5_bF_buf0_), .C(_7630_), .D(_7632__bF_buf3), .Y(_7633_) );
INVX1 INVX1_640 ( .A(_7633_), .Y(_7634_) );
AOI22X1 AOI22X1_48 ( .A(_4584_), .B(_7618_), .C(_7634_), .D(_7622_), .Y(_7635_) );
OAI21X1 OAI21X1_1231 ( .A(_4538__bF_buf0), .B(_7614_), .C(_7635_), .Y(_7636_) );
NAND2X1 NAND2X1_466 ( .A(resetn_bF_buf3), .B(_7636_), .Y(_7637_) );
OAI21X1 OAI21X1_1232 ( .A(_4454_), .B(mem_do_wdata), .C(cpu_state_5_bF_buf3_), .Y(_7638_) );
OAI21X1 OAI21X1_1233 ( .A(_4582_), .B(_4575__bF_buf3), .C(_7627_), .Y(_7639_) );
INVX1 INVX1_641 ( .A(_7639_), .Y(_7640_) );
NAND3X1 NAND3X1_33 ( .A(resetn_bF_buf2), .B(_7638_), .C(_7640_), .Y(_7641_) );
AOI21X1 AOI21X1_315 ( .A(_7630_), .B(_7631__bF_buf4), .C(_7641_), .Y(_7642_) );
OAI21X1 OAI21X1_1234 ( .A(_4491_), .B(_7642_), .C(_7637_), .Y(_81__0_) );
INVX1 INVX1_642 ( .A(_7551__bF_buf2), .Y(_7643_) );
NOR2X1 NOR2X1_508 ( .A(cpuregs_24_[1]), .B(decoded_rs1_0_bF_buf39_), .Y(_7644_) );
OAI21X1 OAI21X1_1235 ( .A(_7569__bF_buf36), .B(cpuregs_25_[1]), .C(_7556__bF_buf32), .Y(_7645_) );
NOR2X1 NOR2X1_509 ( .A(cpuregs_27_[1]), .B(_7569__bF_buf35), .Y(_7646_) );
OAI21X1 OAI21X1_1236 ( .A(cpuregs_26_[1]), .B(decoded_rs1_0_bF_buf38_), .C(decoded_rs1_1_bF_buf32_), .Y(_7647_) );
OAI22X1 OAI22X1_95 ( .A(_7646_), .B(_7647_), .C(_7645_), .D(_7644_), .Y(_7648_) );
NOR2X1 NOR2X1_510 ( .A(decoded_rs1_2_bF_buf6_), .B(_7648_), .Y(_7649_) );
NOR2X1 NOR2X1_511 ( .A(cpuregs_28_[1]), .B(decoded_rs1_0_bF_buf37_), .Y(_7650_) );
OAI21X1 OAI21X1_1237 ( .A(_7569__bF_buf34), .B(cpuregs_29_[1]), .C(_7556__bF_buf31), .Y(_7651_) );
NOR2X1 NOR2X1_512 ( .A(cpuregs_31_[1]), .B(_7569__bF_buf33), .Y(_7652_) );
OAI21X1 OAI21X1_1238 ( .A(cpuregs_30_[1]), .B(decoded_rs1_0_bF_buf36_), .C(decoded_rs1_1_bF_buf31_), .Y(_7653_) );
OAI22X1 OAI22X1_96 ( .A(_7652_), .B(_7653_), .C(_7651_), .D(_7650_), .Y(_7654_) );
OAI21X1 OAI21X1_1239 ( .A(_7654_), .B(_7560__bF_buf8), .C(decoded_rs1_3_bF_buf4_), .Y(_7655_) );
NOR2X1 NOR2X1_513 ( .A(cpuregs_16_[1]), .B(decoded_rs1_0_bF_buf35_), .Y(_7656_) );
OAI21X1 OAI21X1_1240 ( .A(_7569__bF_buf32), .B(cpuregs_17_[1]), .C(_7556__bF_buf30), .Y(_7657_) );
NOR2X1 NOR2X1_514 ( .A(cpuregs_19_[1]), .B(_7569__bF_buf31), .Y(_7658_) );
OAI21X1 OAI21X1_1241 ( .A(cpuregs_18_[1]), .B(decoded_rs1_0_bF_buf34_), .C(decoded_rs1_1_bF_buf30_), .Y(_7659_) );
OAI22X1 OAI22X1_97 ( .A(_7658_), .B(_7659_), .C(_7657_), .D(_7656_), .Y(_7660_) );
NOR2X1 NOR2X1_515 ( .A(cpuregs_20_[1]), .B(decoded_rs1_0_bF_buf33_), .Y(_7661_) );
OAI21X1 OAI21X1_1242 ( .A(_7569__bF_buf30), .B(cpuregs_21_[1]), .C(_7556__bF_buf29), .Y(_7662_) );
NOR2X1 NOR2X1_516 ( .A(cpuregs_23_[1]), .B(_7569__bF_buf29), .Y(_7663_) );
OAI21X1 OAI21X1_1243 ( .A(cpuregs_22_[1]), .B(decoded_rs1_0_bF_buf32_), .C(decoded_rs1_1_bF_buf29_), .Y(_7664_) );
OAI22X1 OAI22X1_98 ( .A(_7663_), .B(_7664_), .C(_7662_), .D(_7661_), .Y(_7665_) );
MUX2X1 MUX2X1_144 ( .A(_7665_), .B(_7660_), .S(decoded_rs1_2_bF_buf5_), .Y(_7666_) );
OAI22X1 OAI22X1_99 ( .A(_7655_), .B(_7649_), .C(_7666_), .D(decoded_rs1_3_bF_buf3_), .Y(_7667_) );
NOR2X1 NOR2X1_517 ( .A(_7552__bF_buf4), .B(_7667_), .Y(_7668_) );
INVX1 INVX1_643 ( .A(cpuregs_9_[1]), .Y(_7669_) );
AOI21X1 AOI21X1_316 ( .A(decoded_rs1_0_bF_buf31_), .B(_7669_), .C(decoded_rs1_1_bF_buf28_), .Y(_7670_) );
OAI21X1 OAI21X1_1244 ( .A(cpuregs_8_[1]), .B(decoded_rs1_0_bF_buf30_), .C(_7670_), .Y(_7671_) );
NOR2X1 NOR2X1_518 ( .A(cpuregs_11_[1]), .B(_7569__bF_buf28), .Y(_7672_) );
OAI21X1 OAI21X1_1245 ( .A(cpuregs_10_[1]), .B(decoded_rs1_0_bF_buf29_), .C(decoded_rs1_1_bF_buf27_), .Y(_7673_) );
OAI21X1 OAI21X1_1246 ( .A(_7672_), .B(_7673_), .C(_7671_), .Y(_7674_) );
NOR2X1 NOR2X1_519 ( .A(decoded_rs1_2_bF_buf4_), .B(_7674_), .Y(_7675_) );
NOR2X1 NOR2X1_520 ( .A(cpuregs_12_[1]), .B(decoded_rs1_0_bF_buf28_), .Y(_7676_) );
OAI21X1 OAI21X1_1247 ( .A(_7569__bF_buf27), .B(cpuregs_13_[1]), .C(_7556__bF_buf28), .Y(_7677_) );
AOI21X1 AOI21X1_317 ( .A(_5427_), .B(_7569__bF_buf26), .C(_7556__bF_buf27), .Y(_7678_) );
OAI21X1 OAI21X1_1248 ( .A(cpuregs_15_[1]), .B(_7569__bF_buf25), .C(_7678_), .Y(_7679_) );
OAI21X1 OAI21X1_1249 ( .A(_7676_), .B(_7677_), .C(_7679_), .Y(_7680_) );
OAI21X1 OAI21X1_1250 ( .A(_7680_), .B(_7560__bF_buf7), .C(decoded_rs1_3_bF_buf2_), .Y(_7681_) );
NOR2X1 NOR2X1_521 ( .A(cpuregs_0_[1]), .B(decoded_rs1_0_bF_buf27_), .Y(_7682_) );
OAI21X1 OAI21X1_1251 ( .A(_7569__bF_buf24), .B(cpuregs_1_[1]), .C(_7556__bF_buf26), .Y(_7683_) );
NOR2X1 NOR2X1_522 ( .A(cpuregs_3_[1]), .B(_7569__bF_buf23), .Y(_7684_) );
OAI21X1 OAI21X1_1252 ( .A(cpuregs_2_[1]), .B(decoded_rs1_0_bF_buf26_), .C(decoded_rs1_1_bF_buf26_), .Y(_7685_) );
OAI22X1 OAI22X1_100 ( .A(_7684_), .B(_7685_), .C(_7683_), .D(_7682_), .Y(_7686_) );
NOR2X1 NOR2X1_523 ( .A(cpuregs_4_[1]), .B(decoded_rs1_0_bF_buf25_), .Y(_7687_) );
OAI21X1 OAI21X1_1253 ( .A(_7569__bF_buf22), .B(cpuregs_5_[1]), .C(_7556__bF_buf25), .Y(_7688_) );
NOR2X1 NOR2X1_524 ( .A(cpuregs_7_[1]), .B(_7569__bF_buf21), .Y(_7689_) );
OAI21X1 OAI21X1_1254 ( .A(cpuregs_6_[1]), .B(decoded_rs1_0_bF_buf24_), .C(decoded_rs1_1_bF_buf25_), .Y(_7690_) );
OAI22X1 OAI22X1_101 ( .A(_7689_), .B(_7690_), .C(_7688_), .D(_7687_), .Y(_7691_) );
MUX2X1 MUX2X1_145 ( .A(_7691_), .B(_7686_), .S(decoded_rs1_2_bF_buf3_), .Y(_7692_) );
OAI22X1 OAI22X1_102 ( .A(decoded_rs1_3_bF_buf1_), .B(_7692_), .C(_7681_), .D(_7675_), .Y(_7693_) );
OAI21X1 OAI21X1_1255 ( .A(_7693_), .B(decoded_rs1_4_bF_buf1_), .C(_7587_), .Y(_7694_) );
OAI22X1 OAI22X1_103 ( .A(_4643_), .B(_7643_), .C(_7694_), .D(_7668_), .Y(_7695_) );
AND2X2 AND2X2_50 ( .A(_7695_), .B(cpu_state_2_bF_buf2_), .Y(_7696_) );
INVX1 INVX1_644 ( .A(_4584_), .Y(_7697_) );
INVX1 INVX1_645 ( .A(_7616_), .Y(_7698_) );
NOR2X1 NOR2X1_525 ( .A(_5179_), .B(_7698__bF_buf4), .Y(_7699_) );
NOR2X1 NOR2X1_526 ( .A(instr_slli), .B(instr_sll), .Y(_7700_) );
NOR2X1 NOR2X1_527 ( .A(_4491_), .B(_7700__bF_buf5), .Y(_7701_) );
NOR2X1 NOR2X1_528 ( .A(_7701_), .B(_4580__bF_buf0), .Y(_7702_) );
OAI21X1 OAI21X1_1256 ( .A(_5148_), .B(_7698__bF_buf3), .C(_7702_), .Y(_7703_) );
OAI21X1 OAI21X1_1257 ( .A(_4579__bF_buf2), .B(_7699_), .C(_7703_), .Y(_7704_) );
XOR2X1 XOR2X1_2 ( .A(_10734__1_), .B(decoded_imm_1_), .Y(_7705_) );
XOR2X1 XOR2X1_3 ( .A(_7705_), .B(_7621_), .Y(_7706_) );
NAND2X1 NAND2X1_467 ( .A(_7706_), .B(_7634_), .Y(_7707_) );
OAI21X1 OAI21X1_1258 ( .A(_7697__bF_buf3), .B(_7704_), .C(_7707_), .Y(_7708_) );
OAI21X1 OAI21X1_1259 ( .A(_7708_), .B(_7696_), .C(resetn_bF_buf1), .Y(_7709_) );
OAI21X1 OAI21X1_1260 ( .A(_4490_), .B(_7642_), .C(_7709_), .Y(_81__1_) );
NOR2X1 NOR2X1_529 ( .A(_4644_), .B(_7643_), .Y(_7710_) );
NAND2X1 NAND2X1_468 ( .A(cpuregs_21_[2]), .B(decoded_rs1_0_bF_buf23_), .Y(_7711_) );
OAI21X1 OAI21X1_1261 ( .A(_5549_), .B(decoded_rs1_0_bF_buf22_), .C(_7711_), .Y(_7712_) );
NAND2X1 NAND2X1_469 ( .A(cpuregs_23_[2]), .B(decoded_rs1_0_bF_buf21_), .Y(_7713_) );
OAI21X1 OAI21X1_1262 ( .A(_5552_), .B(decoded_rs1_0_bF_buf20_), .C(_7713_), .Y(_7714_) );
MUX2X1 MUX2X1_146 ( .A(_7714_), .B(_7712_), .S(decoded_rs1_1_bF_buf24_), .Y(_7715_) );
NAND2X1 NAND2X1_470 ( .A(cpuregs_17_[2]), .B(decoded_rs1_0_bF_buf19_), .Y(_7716_) );
OAI21X1 OAI21X1_1263 ( .A(_5541_), .B(decoded_rs1_0_bF_buf18_), .C(_7716_), .Y(_7717_) );
NAND2X1 NAND2X1_471 ( .A(cpuregs_19_[2]), .B(decoded_rs1_0_bF_buf17_), .Y(_7718_) );
OAI21X1 OAI21X1_1264 ( .A(_5544_), .B(decoded_rs1_0_bF_buf16_), .C(_7718_), .Y(_7719_) );
MUX2X1 MUX2X1_147 ( .A(_7719_), .B(_7717_), .S(decoded_rs1_1_bF_buf23_), .Y(_7720_) );
MUX2X1 MUX2X1_148 ( .A(_7720_), .B(_7715_), .S(_7560__bF_buf6), .Y(_7721_) );
OAI21X1 OAI21X1_1265 ( .A(_5527_), .B(decoded_rs1_0_bF_buf15_), .C(decoded_rs1_1_bF_buf22_), .Y(_7722_) );
AOI21X1 AOI21X1_318 ( .A(cpuregs_27_[2]), .B(decoded_rs1_0_bF_buf14_), .C(_7722_), .Y(_7723_) );
AND2X2 AND2X2_51 ( .A(cpuregs_25_[2]), .B(decoded_rs1_0_bF_buf13_), .Y(_7724_) );
OAI21X1 OAI21X1_1266 ( .A(_5535_), .B(decoded_rs1_0_bF_buf12_), .C(_7556__bF_buf24), .Y(_7725_) );
OAI21X1 OAI21X1_1267 ( .A(_7725_), .B(_7724_), .C(_7560__bF_buf5), .Y(_7726_) );
OAI21X1 OAI21X1_1268 ( .A(_5529_), .B(decoded_rs1_0_bF_buf11_), .C(decoded_rs1_1_bF_buf21_), .Y(_7727_) );
AOI21X1 AOI21X1_319 ( .A(cpuregs_31_[2]), .B(decoded_rs1_0_bF_buf10_), .C(_7727_), .Y(_7728_) );
NOR2X1 NOR2X1_530 ( .A(decoded_rs1_0_bF_buf9_), .B(_5537_), .Y(_7729_) );
OAI21X1 OAI21X1_1269 ( .A(_5532_), .B(_7569__bF_buf20), .C(_7556__bF_buf23), .Y(_7730_) );
OAI21X1 OAI21X1_1270 ( .A(_7730_), .B(_7729_), .C(decoded_rs1_2_bF_buf2_), .Y(_7731_) );
OAI22X1 OAI22X1_104 ( .A(_7726_), .B(_7723_), .C(_7731_), .D(_7728_), .Y(_7732_) );
MUX2X1 MUX2X1_149 ( .A(_7732_), .B(_7721_), .S(decoded_rs1_3_bF_buf0_), .Y(_7733_) );
NOR2X1 NOR2X1_531 ( .A(cpuregs_0_[2]), .B(decoded_rs1_0_bF_buf8_), .Y(_7734_) );
OAI21X1 OAI21X1_1271 ( .A(_7569__bF_buf19), .B(cpuregs_1_[2]), .C(_7556__bF_buf22), .Y(_7735_) );
NOR2X1 NOR2X1_532 ( .A(cpuregs_3_[2]), .B(_7569__bF_buf18), .Y(_7736_) );
OAI21X1 OAI21X1_1272 ( .A(cpuregs_2_[2]), .B(decoded_rs1_0_bF_buf7_), .C(decoded_rs1_1_bF_buf20_), .Y(_7737_) );
OAI22X1 OAI22X1_105 ( .A(_7736_), .B(_7737_), .C(_7735_), .D(_7734_), .Y(_7738_) );
NOR2X1 NOR2X1_533 ( .A(decoded_rs1_2_bF_buf1_), .B(_7738_), .Y(_7739_) );
NOR2X1 NOR2X1_534 ( .A(cpuregs_4_[2]), .B(decoded_rs1_0_bF_buf6_), .Y(_7740_) );
OAI21X1 OAI21X1_1273 ( .A(_7569__bF_buf17), .B(cpuregs_5_[2]), .C(_7556__bF_buf21), .Y(_7741_) );
NOR2X1 NOR2X1_535 ( .A(cpuregs_7_[2]), .B(_7569__bF_buf16), .Y(_7742_) );
OAI21X1 OAI21X1_1274 ( .A(cpuregs_6_[2]), .B(decoded_rs1_0_bF_buf5_), .C(decoded_rs1_1_bF_buf19_), .Y(_7743_) );
OAI22X1 OAI22X1_106 ( .A(_7742_), .B(_7743_), .C(_7741_), .D(_7740_), .Y(_7744_) );
OAI21X1 OAI21X1_1275 ( .A(_7744_), .B(_7560__bF_buf4), .C(_7561__bF_buf2), .Y(_7745_) );
NOR2X1 NOR2X1_536 ( .A(cpuregs_12_[2]), .B(decoded_rs1_0_bF_buf4_), .Y(_7746_) );
OAI21X1 OAI21X1_1276 ( .A(_7569__bF_buf15), .B(cpuregs_13_[2]), .C(_7556__bF_buf20), .Y(_7747_) );
NOR2X1 NOR2X1_537 ( .A(cpuregs_15_[2]), .B(_7569__bF_buf14), .Y(_7748_) );
OAI21X1 OAI21X1_1277 ( .A(cpuregs_14_[2]), .B(decoded_rs1_0_bF_buf3_), .C(decoded_rs1_1_bF_buf18_), .Y(_7749_) );
OAI22X1 OAI22X1_107 ( .A(_7748_), .B(_7749_), .C(_7747_), .D(_7746_), .Y(_7750_) );
NOR2X1 NOR2X1_538 ( .A(_7560__bF_buf3), .B(_7750_), .Y(_7751_) );
NOR2X1 NOR2X1_539 ( .A(cpuregs_8_[2]), .B(decoded_rs1_0_bF_buf2_), .Y(_7752_) );
OAI21X1 OAI21X1_1278 ( .A(_7569__bF_buf13), .B(cpuregs_9_[2]), .C(_7556__bF_buf19), .Y(_7753_) );
NOR2X1 NOR2X1_540 ( .A(cpuregs_11_[2]), .B(_7569__bF_buf12), .Y(_7754_) );
OAI21X1 OAI21X1_1279 ( .A(cpuregs_10_[2]), .B(decoded_rs1_0_bF_buf1_), .C(decoded_rs1_1_bF_buf17_), .Y(_7755_) );
OAI22X1 OAI22X1_108 ( .A(_7754_), .B(_7755_), .C(_7753_), .D(_7752_), .Y(_7756_) );
OAI21X1 OAI21X1_1280 ( .A(_7756_), .B(decoded_rs1_2_bF_buf0_), .C(decoded_rs1_3_bF_buf6_), .Y(_7757_) );
OAI22X1 OAI22X1_109 ( .A(_7745_), .B(_7739_), .C(_7751_), .D(_7757_), .Y(_7758_) );
OAI21X1 OAI21X1_1281 ( .A(_7758_), .B(decoded_rs1_4_bF_buf0_), .C(_7587_), .Y(_7759_) );
AOI21X1 AOI21X1_320 ( .A(decoded_rs1_4_bF_buf4_), .B(_7733_), .C(_7759_), .Y(_7760_) );
OAI21X1 OAI21X1_1282 ( .A(_7760_), .B(_7710_), .C(cpu_state_2_bF_buf1_), .Y(_7761_) );
INVX1 INVX1_646 ( .A(decoded_imm_1_), .Y(_7762_) );
NAND2X1 NAND2X1_472 ( .A(_7621_), .B(_7705_), .Y(_7763_) );
OAI21X1 OAI21X1_1283 ( .A(_4490_), .B(_7762_), .C(_7763_), .Y(_7764_) );
NAND2X1 NAND2X1_473 ( .A(_10734__2_), .B(decoded_imm_2_), .Y(_7765_) );
INVX1 INVX1_647 ( .A(decoded_imm_2_), .Y(_7766_) );
NAND2X1 NAND2X1_474 ( .A(_5148_), .B(_7766_), .Y(_7767_) );
NAND2X1 NAND2X1_475 ( .A(_7765_), .B(_7767_), .Y(_7768_) );
XNOR2X1 XNOR2X1_2 ( .A(_7764_), .B(_7768_), .Y(_7769_) );
NOR2X1 NOR2X1_541 ( .A(_7623__bF_buf3), .B(_7769_), .Y(_7770_) );
OAI21X1 OAI21X1_1284 ( .A(_7624__bF_buf3), .B(_10734__2_), .C(cpu_state_5_bF_buf2_), .Y(_7771_) );
INVX1 INVX1_648 ( .A(_7769_), .Y(_7772_) );
OAI21X1 OAI21X1_1285 ( .A(_4454_), .B(mem_do_rdata), .C(_10734__2_), .Y(_7773_) );
OAI21X1 OAI21X1_1286 ( .A(_7772_), .B(_7631__bF_buf3), .C(_7773_), .Y(_7774_) );
NOR2X1 NOR2X1_542 ( .A(_4490_), .B(_7700__bF_buf4), .Y(_7775_) );
AOI21X1 AOI21X1_321 ( .A(_10734__3_), .B(_7616_), .C(_7775_), .Y(_7776_) );
NOR2X1 NOR2X1_543 ( .A(_7776_), .B(_4580__bF_buf4), .Y(_7777_) );
INVX1 INVX1_649 ( .A(_7615_), .Y(_7778_) );
OAI21X1 OAI21X1_1287 ( .A(_7778_), .B(_7700__bF_buf3), .C(_10734__6_), .Y(_7779_) );
NOR2X1 NOR2X1_544 ( .A(_4579__bF_buf1), .B(_7779_), .Y(_7780_) );
OAI21X1 OAI21X1_1288 ( .A(_7777_), .B(_7780_), .C(_4584_), .Y(_7781_) );
OAI21X1 OAI21X1_1289 ( .A(_5148_), .B(_7640_), .C(_7781_), .Y(_7782_) );
AOI21X1 AOI21X1_322 ( .A(_7630_), .B(_7774_), .C(_7782_), .Y(_7783_) );
OAI21X1 OAI21X1_1290 ( .A(_7770_), .B(_7771_), .C(_7783_), .Y(_7784_) );
NOR2X1 NOR2X1_545 ( .A(_4426__bF_buf11), .B(_7784_), .Y(_7785_) );
AOI22X1 AOI22X1_49 ( .A(_4426__bF_buf10), .B(_5148_), .C(_7785_), .D(_7761_), .Y(_81__2_) );
INVX1 INVX1_650 ( .A(reg_pc_3_), .Y(_7786_) );
AOI21X1 AOI21X1_323 ( .A(decoded_rs1_1_bF_buf16_), .B(_5614_), .C(decoded_rs1_0_bF_buf0_), .Y(_7787_) );
OAI21X1 OAI21X1_1291 ( .A(cpuregs_16_[3]), .B(decoded_rs1_1_bF_buf15_), .C(_7787_), .Y(_7788_) );
NOR2X1 NOR2X1_546 ( .A(cpuregs_17_[3]), .B(decoded_rs1_1_bF_buf14_), .Y(_7789_) );
OAI21X1 OAI21X1_1292 ( .A(_7556__bF_buf18), .B(cpuregs_19_[3]), .C(decoded_rs1_0_bF_buf57_), .Y(_7790_) );
OAI21X1 OAI21X1_1293 ( .A(_7789_), .B(_7790_), .C(_7788_), .Y(_7791_) );
NOR2X1 NOR2X1_547 ( .A(decoded_rs1_2_bF_buf12_), .B(_7791_), .Y(_7792_) );
NOR2X1 NOR2X1_548 ( .A(cpuregs_20_[3]), .B(decoded_rs1_1_bF_buf13_), .Y(_7793_) );
OAI21X1 OAI21X1_1294 ( .A(_7556__bF_buf17), .B(cpuregs_22_[3]), .C(_7569__bF_buf11), .Y(_7794_) );
AOI21X1 AOI21X1_324 ( .A(decoded_rs1_1_bF_buf12_), .B(_5621_), .C(_7569__bF_buf10), .Y(_7795_) );
OAI21X1 OAI21X1_1295 ( .A(cpuregs_21_[3]), .B(decoded_rs1_1_bF_buf11_), .C(_7795_), .Y(_7796_) );
OAI21X1 OAI21X1_1296 ( .A(_7793_), .B(_7794_), .C(_7796_), .Y(_7797_) );
OAI21X1 OAI21X1_1297 ( .A(_7797_), .B(_7560__bF_buf2), .C(_7561__bF_buf1), .Y(_7798_) );
NOR2X1 NOR2X1_549 ( .A(cpuregs_24_[3]), .B(decoded_rs1_0_bF_buf56_), .Y(_7799_) );
OAI21X1 OAI21X1_1298 ( .A(_7569__bF_buf9), .B(cpuregs_25_[3]), .C(_7556__bF_buf16), .Y(_7800_) );
NOR2X1 NOR2X1_550 ( .A(cpuregs_27_[3]), .B(_7569__bF_buf8), .Y(_7801_) );
OAI21X1 OAI21X1_1299 ( .A(cpuregs_26_[3]), .B(decoded_rs1_0_bF_buf55_), .C(decoded_rs1_1_bF_buf10_), .Y(_7802_) );
OAI22X1 OAI22X1_110 ( .A(_7801_), .B(_7802_), .C(_7800_), .D(_7799_), .Y(_7803_) );
NOR2X1 NOR2X1_551 ( .A(decoded_rs1_2_bF_buf11_), .B(_7803_), .Y(_7804_) );
NOR2X1 NOR2X1_552 ( .A(cpuregs_28_[3]), .B(decoded_rs1_0_bF_buf54_), .Y(_7805_) );
OAI21X1 OAI21X1_1300 ( .A(_7569__bF_buf7), .B(cpuregs_29_[3]), .C(_7556__bF_buf15), .Y(_7806_) );
NOR2X1 NOR2X1_553 ( .A(cpuregs_31_[3]), .B(_7569__bF_buf6), .Y(_7807_) );
OAI21X1 OAI21X1_1301 ( .A(cpuregs_30_[3]), .B(decoded_rs1_0_bF_buf53_), .C(decoded_rs1_1_bF_buf9_), .Y(_7808_) );
OAI22X1 OAI22X1_111 ( .A(_7807_), .B(_7808_), .C(_7806_), .D(_7805_), .Y(_7809_) );
OAI21X1 OAI21X1_1302 ( .A(_7809_), .B(_7560__bF_buf1), .C(decoded_rs1_3_bF_buf5_), .Y(_7810_) );
OAI22X1 OAI22X1_112 ( .A(_7804_), .B(_7810_), .C(_7798_), .D(_7792_), .Y(_7811_) );
NOR2X1 NOR2X1_554 ( .A(_7552__bF_buf3), .B(_7811_), .Y(_7812_) );
NOR2X1 NOR2X1_555 ( .A(cpuregs_0_[3]), .B(decoded_rs1_0_bF_buf52_), .Y(_7813_) );
OAI21X1 OAI21X1_1303 ( .A(_7569__bF_buf5), .B(cpuregs_1_[3]), .C(_7556__bF_buf14), .Y(_7814_) );
NOR2X1 NOR2X1_556 ( .A(cpuregs_3_[3]), .B(_7569__bF_buf4), .Y(_7815_) );
OAI21X1 OAI21X1_1304 ( .A(cpuregs_2_[3]), .B(decoded_rs1_0_bF_buf51_), .C(decoded_rs1_1_bF_buf8_), .Y(_7816_) );
OAI22X1 OAI22X1_113 ( .A(_7815_), .B(_7816_), .C(_7814_), .D(_7813_), .Y(_7817_) );
NOR2X1 NOR2X1_557 ( .A(decoded_rs1_2_bF_buf10_), .B(_7817_), .Y(_7818_) );
NOR2X1 NOR2X1_558 ( .A(cpuregs_4_[3]), .B(decoded_rs1_0_bF_buf50_), .Y(_7819_) );
OAI21X1 OAI21X1_1305 ( .A(_7569__bF_buf3), .B(cpuregs_5_[3]), .C(_7556__bF_buf13), .Y(_7820_) );
NOR2X1 NOR2X1_559 ( .A(cpuregs_7_[3]), .B(_7569__bF_buf2), .Y(_7821_) );
OAI21X1 OAI21X1_1306 ( .A(cpuregs_6_[3]), .B(decoded_rs1_0_bF_buf49_), .C(decoded_rs1_1_bF_buf7_), .Y(_7822_) );
OAI22X1 OAI22X1_114 ( .A(_7821_), .B(_7822_), .C(_7820_), .D(_7819_), .Y(_7823_) );
OAI21X1 OAI21X1_1307 ( .A(_7823_), .B(_7560__bF_buf0), .C(_7561__bF_buf0), .Y(_7824_) );
NOR2X1 NOR2X1_560 ( .A(cpuregs_12_[3]), .B(decoded_rs1_0_bF_buf48_), .Y(_7825_) );
OAI21X1 OAI21X1_1308 ( .A(_7569__bF_buf1), .B(cpuregs_13_[3]), .C(_7556__bF_buf12), .Y(_7826_) );
NOR2X1 NOR2X1_561 ( .A(cpuregs_15_[3]), .B(_7569__bF_buf0), .Y(_7827_) );
OAI21X1 OAI21X1_1309 ( .A(cpuregs_14_[3]), .B(decoded_rs1_0_bF_buf47_), .C(decoded_rs1_1_bF_buf6_), .Y(_7828_) );
OAI22X1 OAI22X1_115 ( .A(_7827_), .B(_7828_), .C(_7826_), .D(_7825_), .Y(_7829_) );
NOR2X1 NOR2X1_562 ( .A(_7560__bF_buf12), .B(_7829_), .Y(_7830_) );
NOR2X1 NOR2X1_563 ( .A(cpuregs_8_[3]), .B(decoded_rs1_0_bF_buf46_), .Y(_7831_) );
OAI21X1 OAI21X1_1310 ( .A(_7569__bF_buf48), .B(cpuregs_9_[3]), .C(_7556__bF_buf11), .Y(_7832_) );
NOR2X1 NOR2X1_564 ( .A(cpuregs_11_[3]), .B(_7569__bF_buf47), .Y(_7833_) );
OAI21X1 OAI21X1_1311 ( .A(cpuregs_10_[3]), .B(decoded_rs1_0_bF_buf45_), .C(decoded_rs1_1_bF_buf5_), .Y(_7834_) );
OAI22X1 OAI22X1_116 ( .A(_7833_), .B(_7834_), .C(_7832_), .D(_7831_), .Y(_7835_) );
OAI21X1 OAI21X1_1312 ( .A(_7835_), .B(decoded_rs1_2_bF_buf9_), .C(decoded_rs1_3_bF_buf4_), .Y(_7836_) );
OAI22X1 OAI22X1_117 ( .A(_7824_), .B(_7818_), .C(_7830_), .D(_7836_), .Y(_7837_) );
OAI21X1 OAI21X1_1313 ( .A(_7837_), .B(decoded_rs1_4_bF_buf3_), .C(_7587_), .Y(_7838_) );
OAI22X1 OAI22X1_118 ( .A(_7786_), .B(_7643_), .C(_7812_), .D(_7838_), .Y(_7839_) );
AND2X2 AND2X2_52 ( .A(_7839_), .B(cpu_state_2_bF_buf0_), .Y(_7840_) );
NOR2X1 NOR2X1_565 ( .A(_5148_), .B(_7700__bF_buf2), .Y(_7841_) );
AOI21X1 AOI21X1_325 ( .A(_10734__4_), .B(_7616_), .C(_7841_), .Y(_7842_) );
NOR2X1 NOR2X1_566 ( .A(_7842_), .B(_4580__bF_buf3), .Y(_7843_) );
OAI21X1 OAI21X1_1314 ( .A(_7778_), .B(_7700__bF_buf1), .C(_10734__7_), .Y(_7844_) );
NOR2X1 NOR2X1_567 ( .A(_4579__bF_buf0), .B(_7844_), .Y(_7845_) );
OAI21X1 OAI21X1_1315 ( .A(_7843_), .B(_7845_), .C(_4584_), .Y(_7846_) );
INVX1 INVX1_651 ( .A(_7765_), .Y(_7847_) );
AOI21X1 AOI21X1_326 ( .A(_7767_), .B(_7764_), .C(_7847_), .Y(_7848_) );
NAND2X1 NAND2X1_476 ( .A(_10734__3_), .B(decoded_imm_3_), .Y(_7849_) );
INVX1 INVX1_652 ( .A(decoded_imm_3_), .Y(_7850_) );
NAND2X1 NAND2X1_477 ( .A(_5130_), .B(_7850_), .Y(_7851_) );
NAND2X1 NAND2X1_478 ( .A(_7849_), .B(_7851_), .Y(_7852_) );
XNOR2X1 XNOR2X1_3 ( .A(_7848_), .B(_7852_), .Y(_7853_) );
OAI21X1 OAI21X1_1316 ( .A(_7633_), .B(_7853_), .C(_7846_), .Y(_7854_) );
OAI21X1 OAI21X1_1317 ( .A(_7840_), .B(_7854_), .C(resetn_bF_buf0), .Y(_7855_) );
OAI21X1 OAI21X1_1318 ( .A(_5130_), .B(_7642_), .C(_7855_), .Y(_81__3_) );
AOI21X1 AOI21X1_327 ( .A(cpuregs_26_[4]), .B(_7569__bF_buf46), .C(_7556__bF_buf10), .Y(_7856_) );
OAI21X1 OAI21X1_1319 ( .A(_5670_), .B(_7569__bF_buf45), .C(_7856_), .Y(_7857_) );
OAI21X1 OAI21X1_1320 ( .A(_5667_), .B(decoded_rs1_0_bF_buf44_), .C(_7556__bF_buf9), .Y(_7858_) );
AOI21X1 AOI21X1_328 ( .A(cpuregs_25_[4]), .B(decoded_rs1_0_bF_buf43_), .C(_7858_), .Y(_7859_) );
NOR2X1 NOR2X1_568 ( .A(decoded_rs1_2_bF_buf8_), .B(_7859_), .Y(_7860_) );
NOR2X1 NOR2X1_569 ( .A(cpuregs_28_[4]), .B(decoded_rs1_0_bF_buf42_), .Y(_7861_) );
OAI21X1 OAI21X1_1321 ( .A(_7569__bF_buf44), .B(cpuregs_29_[4]), .C(_7556__bF_buf8), .Y(_7862_) );
NOR2X1 NOR2X1_570 ( .A(cpuregs_31_[4]), .B(_7569__bF_buf43), .Y(_7863_) );
OAI21X1 OAI21X1_1322 ( .A(cpuregs_30_[4]), .B(decoded_rs1_0_bF_buf41_), .C(decoded_rs1_1_bF_buf4_), .Y(_7864_) );
OAI22X1 OAI22X1_119 ( .A(_7863_), .B(_7864_), .C(_7862_), .D(_7861_), .Y(_7865_) );
AOI22X1 AOI22X1_50 ( .A(decoded_rs1_2_bF_buf7_), .B(_7865_), .C(_7860_), .D(_7857_), .Y(_7866_) );
AOI21X1 AOI21X1_329 ( .A(decoded_rs1_1_bF_buf3_), .B(_5685_), .C(decoded_rs1_0_bF_buf40_), .Y(_7867_) );
OAI21X1 OAI21X1_1323 ( .A(cpuregs_16_[4]), .B(decoded_rs1_1_bF_buf2_), .C(_7867_), .Y(_7868_) );
NOR2X1 NOR2X1_571 ( .A(cpuregs_17_[4]), .B(decoded_rs1_1_bF_buf1_), .Y(_7869_) );
OAI21X1 OAI21X1_1324 ( .A(_7556__bF_buf7), .B(cpuregs_19_[4]), .C(decoded_rs1_0_bF_buf39_), .Y(_7870_) );
OAI21X1 OAI21X1_1325 ( .A(_7869_), .B(_7870_), .C(_7868_), .Y(_7871_) );
NOR2X1 NOR2X1_572 ( .A(decoded_rs1_2_bF_buf6_), .B(_7871_), .Y(_7872_) );
NOR2X1 NOR2X1_573 ( .A(cpuregs_20_[4]), .B(decoded_rs1_1_bF_buf0_), .Y(_7873_) );
OAI21X1 OAI21X1_1326 ( .A(_7556__bF_buf6), .B(cpuregs_22_[4]), .C(_7569__bF_buf42), .Y(_7874_) );
AOI21X1 AOI21X1_330 ( .A(decoded_rs1_1_bF_buf44_), .B(_5692_), .C(_7569__bF_buf41), .Y(_7875_) );
OAI21X1 OAI21X1_1327 ( .A(cpuregs_21_[4]), .B(decoded_rs1_1_bF_buf43_), .C(_7875_), .Y(_7876_) );
OAI21X1 OAI21X1_1328 ( .A(_7873_), .B(_7874_), .C(_7876_), .Y(_7877_) );
OAI21X1 OAI21X1_1329 ( .A(_7877_), .B(_7560__bF_buf11), .C(_7561__bF_buf6), .Y(_7878_) );
OAI22X1 OAI22X1_120 ( .A(_7878_), .B(_7872_), .C(_7866_), .D(_7561__bF_buf5), .Y(_7879_) );
NOR2X1 NOR2X1_574 ( .A(_7552__bF_buf2), .B(_7879_), .Y(_7880_) );
NOR2X1 NOR2X1_575 ( .A(cpuregs_0_[4]), .B(decoded_rs1_0_bF_buf38_), .Y(_7881_) );
OAI21X1 OAI21X1_1330 ( .A(_7569__bF_buf40), .B(cpuregs_1_[4]), .C(_7556__bF_buf5), .Y(_7882_) );
NOR2X1 NOR2X1_576 ( .A(cpuregs_3_[4]), .B(_7569__bF_buf39), .Y(_7883_) );
OAI21X1 OAI21X1_1331 ( .A(cpuregs_2_[4]), .B(decoded_rs1_0_bF_buf37_), .C(decoded_rs1_1_bF_buf42_), .Y(_7884_) );
OAI22X1 OAI22X1_121 ( .A(_7883_), .B(_7884_), .C(_7882_), .D(_7881_), .Y(_7885_) );
NOR2X1 NOR2X1_577 ( .A(decoded_rs1_2_bF_buf5_), .B(_7885_), .Y(_7886_) );
NOR2X1 NOR2X1_578 ( .A(cpuregs_4_[4]), .B(decoded_rs1_0_bF_buf36_), .Y(_7887_) );
OAI21X1 OAI21X1_1332 ( .A(_7569__bF_buf38), .B(cpuregs_5_[4]), .C(_7556__bF_buf4), .Y(_7888_) );
NOR2X1 NOR2X1_579 ( .A(cpuregs_7_[4]), .B(_7569__bF_buf37), .Y(_7889_) );
OAI21X1 OAI21X1_1333 ( .A(cpuregs_6_[4]), .B(decoded_rs1_0_bF_buf35_), .C(decoded_rs1_1_bF_buf41_), .Y(_7890_) );
OAI22X1 OAI22X1_122 ( .A(_7889_), .B(_7890_), .C(_7888_), .D(_7887_), .Y(_7891_) );
OAI21X1 OAI21X1_1334 ( .A(_7891_), .B(_7560__bF_buf10), .C(_7561__bF_buf4), .Y(_7892_) );
NOR2X1 NOR2X1_580 ( .A(cpuregs_12_[4]), .B(decoded_rs1_0_bF_buf34_), .Y(_7893_) );
OAI21X1 OAI21X1_1335 ( .A(_7569__bF_buf36), .B(cpuregs_13_[4]), .C(_7556__bF_buf3), .Y(_7894_) );
NOR2X1 NOR2X1_581 ( .A(cpuregs_15_[4]), .B(_7569__bF_buf35), .Y(_7895_) );
OAI21X1 OAI21X1_1336 ( .A(cpuregs_14_[4]), .B(decoded_rs1_0_bF_buf33_), .C(decoded_rs1_1_bF_buf40_), .Y(_7896_) );
OAI22X1 OAI22X1_123 ( .A(_7895_), .B(_7896_), .C(_7894_), .D(_7893_), .Y(_7897_) );
NOR2X1 NOR2X1_582 ( .A(_7560__bF_buf9), .B(_7897_), .Y(_7898_) );
NOR2X1 NOR2X1_583 ( .A(cpuregs_8_[4]), .B(decoded_rs1_0_bF_buf32_), .Y(_7899_) );
OAI21X1 OAI21X1_1337 ( .A(_7569__bF_buf34), .B(cpuregs_9_[4]), .C(_7556__bF_buf2), .Y(_7900_) );
NOR2X1 NOR2X1_584 ( .A(cpuregs_11_[4]), .B(_7569__bF_buf33), .Y(_7901_) );
OAI21X1 OAI21X1_1338 ( .A(cpuregs_10_[4]), .B(decoded_rs1_0_bF_buf31_), .C(decoded_rs1_1_bF_buf39_), .Y(_7902_) );
OAI22X1 OAI22X1_124 ( .A(_7901_), .B(_7902_), .C(_7900_), .D(_7899_), .Y(_7903_) );
OAI21X1 OAI21X1_1339 ( .A(_7903_), .B(decoded_rs1_2_bF_buf4_), .C(decoded_rs1_3_bF_buf3_), .Y(_7904_) );
OAI22X1 OAI22X1_125 ( .A(_7892_), .B(_7886_), .C(_7898_), .D(_7904_), .Y(_7905_) );
OAI21X1 OAI21X1_1340 ( .A(_7905_), .B(decoded_rs1_4_bF_buf2_), .C(_7587_), .Y(_7906_) );
OAI22X1 OAI22X1_126 ( .A(_4642_), .B(_7643_), .C(_7880_), .D(_7906_), .Y(_7907_) );
NOR2X1 NOR2X1_585 ( .A(_5130_), .B(_7700__bF_buf0), .Y(_7908_) );
OAI21X1 OAI21X1_1341 ( .A(_7699_), .B(_7908_), .C(_4579__bF_buf4), .Y(_7909_) );
AOI21X1 AOI21X1_331 ( .A(_10734__8_), .B(_7616_), .C(_7701_), .Y(_7910_) );
OAI21X1 OAI21X1_1342 ( .A(_4579__bF_buf3), .B(_7910_), .C(_7909_), .Y(_7911_) );
NAND2X1 NAND2X1_479 ( .A(_7911_), .B(_4584_), .Y(_7912_) );
NOR2X1 NOR2X1_586 ( .A(_10734__4_), .B(decoded_imm_4_), .Y(_7913_) );
INVX1 INVX1_653 ( .A(decoded_imm_4_), .Y(_7914_) );
NOR2X1 NOR2X1_587 ( .A(_5180_), .B(_7914_), .Y(_7915_) );
NOR2X1 NOR2X1_588 ( .A(_7913_), .B(_7915_), .Y(_7916_) );
OAI21X1 OAI21X1_1343 ( .A(_7852_), .B(_7765_), .C(_7849_), .Y(_7917_) );
NOR2X1 NOR2X1_589 ( .A(_7768_), .B(_7852_), .Y(_7918_) );
AOI21X1 AOI21X1_332 ( .A(_7918_), .B(_7764_), .C(_7917_), .Y(_7919_) );
XOR2X1 XOR2X1_4 ( .A(_7919_), .B(_7916_), .Y(_7920_) );
OAI21X1 OAI21X1_1344 ( .A(_7633_), .B(_7920_), .C(_7912_), .Y(_7921_) );
AOI21X1 AOI21X1_333 ( .A(cpu_state_2_bF_buf5_), .B(_7907_), .C(_7921_), .Y(_7922_) );
OAI22X1 OAI22X1_127 ( .A(_5180_), .B(_7642_), .C(_7922_), .D(_4426__bF_buf9), .Y(_81__4_) );
NAND2X1 NAND2X1_480 ( .A(_10734__4_), .B(decoded_imm_4_), .Y(_7923_) );
OAI21X1 OAI21X1_1345 ( .A(_7919_), .B(_7913_), .C(_7923_), .Y(_7924_) );
NAND2X1 NAND2X1_481 ( .A(_10734__5_), .B(decoded_imm_5_), .Y(_7925_) );
INVX1 INVX1_654 ( .A(decoded_imm_5_), .Y(_7926_) );
NAND2X1 NAND2X1_482 ( .A(_5179_), .B(_7926_), .Y(_7927_) );
NAND2X1 NAND2X1_483 ( .A(_7925_), .B(_7927_), .Y(_7928_) );
XNOR2X1 XNOR2X1_4 ( .A(_7924_), .B(_7928_), .Y(_7929_) );
AOI21X1 AOI21X1_334 ( .A(_5179_), .B(_7631__bF_buf2), .C(_7629__bF_buf2), .Y(_7930_) );
OAI21X1 OAI21X1_1346 ( .A(_7929_), .B(_7631__bF_buf1), .C(_7930_), .Y(_7931_) );
AOI21X1 AOI21X1_335 ( .A(_5179_), .B(_7623__bF_buf2), .C(_4587__bF_buf2), .Y(_7932_) );
OAI21X1 OAI21X1_1347 ( .A(_7929_), .B(_7623__bF_buf1), .C(_7932_), .Y(_7933_) );
INVX1 INVX1_655 ( .A(reg_pc_5_), .Y(_7934_) );
NOR2X1 NOR2X1_590 ( .A(cpuregs_1_[5]), .B(decoded_rs1_2_bF_buf3_), .Y(_7935_) );
OAI21X1 OAI21X1_1348 ( .A(_7560__bF_buf8), .B(cpuregs_5_[5]), .C(decoded_rs1_0_bF_buf30_), .Y(_7936_) );
NOR2X1 NOR2X1_591 ( .A(_7935_), .B(_7936_), .Y(_7937_) );
NOR2X1 NOR2X1_592 ( .A(cpuregs_0_[5]), .B(decoded_rs1_2_bF_buf2_), .Y(_7938_) );
OAI21X1 OAI21X1_1349 ( .A(_7560__bF_buf7), .B(cpuregs_4_[5]), .C(_7569__bF_buf32), .Y(_7939_) );
OAI21X1 OAI21X1_1350 ( .A(_7939_), .B(_7938_), .C(_7556__bF_buf1), .Y(_7940_) );
NOR2X1 NOR2X1_593 ( .A(cpuregs_3_[5]), .B(decoded_rs1_2_bF_buf1_), .Y(_7941_) );
OAI21X1 OAI21X1_1351 ( .A(_7560__bF_buf6), .B(cpuregs_7_[5]), .C(decoded_rs1_0_bF_buf29_), .Y(_7942_) );
NOR2X1 NOR2X1_594 ( .A(_7941_), .B(_7942_), .Y(_7943_) );
NOR2X1 NOR2X1_595 ( .A(cpuregs_2_[5]), .B(decoded_rs1_2_bF_buf0_), .Y(_7944_) );
OAI21X1 OAI21X1_1352 ( .A(_7560__bF_buf5), .B(cpuregs_6_[5]), .C(_7569__bF_buf31), .Y(_7945_) );
OAI21X1 OAI21X1_1353 ( .A(_7945_), .B(_7944_), .C(decoded_rs1_1_bF_buf38_), .Y(_7946_) );
OAI22X1 OAI22X1_128 ( .A(_7940_), .B(_7937_), .C(_7943_), .D(_7946_), .Y(_7947_) );
OAI21X1 OAI21X1_1354 ( .A(_5906_), .B(decoded_rs1_0_bF_buf28_), .C(_7556__bF_buf0), .Y(_7948_) );
AOI21X1 AOI21X1_336 ( .A(cpuregs_17_[5]), .B(decoded_rs1_0_bF_buf27_), .C(_7948_), .Y(_7949_) );
INVX1 INVX1_656 ( .A(cpuregs_19_[5]), .Y(_7950_) );
OAI21X1 OAI21X1_1355 ( .A(_7950_), .B(_7569__bF_buf30), .C(decoded_rs1_1_bF_buf37_), .Y(_7951_) );
AOI21X1 AOI21X1_337 ( .A(cpuregs_18_[5]), .B(_7569__bF_buf29), .C(_7951_), .Y(_7952_) );
OAI21X1 OAI21X1_1356 ( .A(_7949_), .B(_7952_), .C(_7560__bF_buf4), .Y(_7953_) );
OAI21X1 OAI21X1_1357 ( .A(_5914_), .B(decoded_rs1_0_bF_buf26_), .C(_7556__bF_buf42), .Y(_7954_) );
AOI21X1 AOI21X1_338 ( .A(cpuregs_21_[5]), .B(decoded_rs1_0_bF_buf25_), .C(_7954_), .Y(_7955_) );
OAI21X1 OAI21X1_1358 ( .A(_5917_), .B(_7569__bF_buf28), .C(decoded_rs1_1_bF_buf36_), .Y(_7956_) );
AOI21X1 AOI21X1_339 ( .A(cpuregs_22_[5]), .B(_7569__bF_buf27), .C(_7956_), .Y(_7957_) );
OAI21X1 OAI21X1_1359 ( .A(_7955_), .B(_7957_), .C(decoded_rs1_2_bF_buf12_), .Y(_7958_) );
AND2X2 AND2X2_53 ( .A(_7953_), .B(_7958_), .Y(_7959_) );
OAI21X1 OAI21X1_1360 ( .A(_7959_), .B(_7552__bF_buf1), .C(_7561__bF_buf3), .Y(_7960_) );
AOI21X1 AOI21X1_340 ( .A(_7552__bF_buf0), .B(_7947_), .C(_7960_), .Y(_7961_) );
OAI21X1 OAI21X1_1361 ( .A(cpuregs_24_[5]), .B(decoded_rs1_1_bF_buf35_), .C(_7569__bF_buf26), .Y(_7962_) );
AOI21X1 AOI21X1_341 ( .A(_5891_), .B(decoded_rs1_1_bF_buf34_), .C(_7962_), .Y(_7963_) );
NOR2X1 NOR2X1_596 ( .A(cpuregs_27_[5]), .B(_7556__bF_buf41), .Y(_7964_) );
OAI21X1 OAI21X1_1362 ( .A(cpuregs_25_[5]), .B(decoded_rs1_1_bF_buf33_), .C(decoded_rs1_0_bF_buf24_), .Y(_7965_) );
NOR2X1 NOR2X1_597 ( .A(_7965_), .B(_7964_), .Y(_7966_) );
OAI21X1 OAI21X1_1363 ( .A(_7963_), .B(_7966_), .C(_7560__bF_buf3), .Y(_7967_) );
AOI21X1 AOI21X1_342 ( .A(_5898_), .B(_7556__bF_buf40), .C(decoded_rs1_0_bF_buf23_), .Y(_7968_) );
OAI21X1 OAI21X1_1364 ( .A(cpuregs_30_[5]), .B(_7556__bF_buf39), .C(_7968_), .Y(_7969_) );
NOR2X1 NOR2X1_598 ( .A(cpuregs_31_[5]), .B(_7556__bF_buf38), .Y(_7970_) );
OAI21X1 OAI21X1_1365 ( .A(cpuregs_29_[5]), .B(decoded_rs1_1_bF_buf32_), .C(decoded_rs1_0_bF_buf22_), .Y(_7971_) );
OAI21X1 OAI21X1_1366 ( .A(_7970_), .B(_7971_), .C(_7969_), .Y(_7972_) );
AOI21X1 AOI21X1_343 ( .A(decoded_rs1_2_bF_buf11_), .B(_7972_), .C(_7552__bF_buf5), .Y(_7973_) );
AOI21X1 AOI21X1_344 ( .A(_4623_), .B(_7556__bF_buf37), .C(decoded_rs1_0_bF_buf21_), .Y(_7974_) );
OAI21X1 OAI21X1_1367 ( .A(cpuregs_10_[5]), .B(_7556__bF_buf36), .C(_7974_), .Y(_7975_) );
AOI21X1 AOI21X1_345 ( .A(_5875_), .B(_7556__bF_buf35), .C(_7569__bF_buf25), .Y(_7976_) );
OAI21X1 OAI21X1_1368 ( .A(cpuregs_11_[5]), .B(_7556__bF_buf34), .C(_7976_), .Y(_7977_) );
AOI21X1 AOI21X1_346 ( .A(_7975_), .B(_7977_), .C(decoded_rs1_2_bF_buf10_), .Y(_7978_) );
AND2X2 AND2X2_54 ( .A(cpuregs_13_[5]), .B(decoded_rs1_0_bF_buf20_), .Y(_7979_) );
INVX1 INVX1_657 ( .A(cpuregs_12_[5]), .Y(_7980_) );
OAI21X1 OAI21X1_1369 ( .A(_7980_), .B(decoded_rs1_0_bF_buf19_), .C(_7556__bF_buf33), .Y(_7981_) );
AOI21X1 AOI21X1_347 ( .A(cpuregs_15_[5]), .B(decoded_rs1_0_bF_buf18_), .C(_7556__bF_buf32), .Y(_7982_) );
OAI21X1 OAI21X1_1370 ( .A(_5884_), .B(decoded_rs1_0_bF_buf17_), .C(_7982_), .Y(_7983_) );
OAI21X1 OAI21X1_1371 ( .A(_7979_), .B(_7981_), .C(_7983_), .Y(_7984_) );
OAI21X1 OAI21X1_1372 ( .A(_7984_), .B(_7560__bF_buf2), .C(_7552__bF_buf4), .Y(_7985_) );
OAI21X1 OAI21X1_1373 ( .A(_7985_), .B(_7978_), .C(decoded_rs1_3_bF_buf2_), .Y(_7986_) );
AOI21X1 AOI21X1_348 ( .A(_7967_), .B(_7973_), .C(_7986_), .Y(_7987_) );
OAI21X1 OAI21X1_1374 ( .A(_7961_), .B(_7987_), .C(_7587_), .Y(_7988_) );
OAI21X1 OAI21X1_1375 ( .A(_7934_), .B(_7643_), .C(_7988_), .Y(_7989_) );
OAI21X1 OAI21X1_1376 ( .A(_7778_), .B(_7700__bF_buf5), .C(_10734__9_), .Y(_7990_) );
NOR2X1 NOR2X1_599 ( .A(_7775_), .B(_4579__bF_buf2), .Y(_7991_) );
NOR2X1 NOR2X1_600 ( .A(_5180_), .B(_7700__bF_buf4), .Y(_7992_) );
NOR2X1 NOR2X1_601 ( .A(_7992_), .B(_4580__bF_buf2), .Y(_7993_) );
AOI22X1 AOI22X1_51 ( .A(_7990_), .B(_7991_), .C(_7993_), .D(_7779_), .Y(_7994_) );
AOI21X1 AOI21X1_349 ( .A(_7994_), .B(_4584_), .C(_4426__bF_buf8), .Y(_7995_) );
OAI21X1 OAI21X1_1377 ( .A(_5179_), .B(_7640_), .C(_7995_), .Y(_7996_) );
AOI21X1 AOI21X1_350 ( .A(cpu_state_2_bF_buf4_), .B(_7989_), .C(_7996_), .Y(_7997_) );
AND2X2 AND2X2_55 ( .A(_7997_), .B(_7933_), .Y(_7998_) );
AOI22X1 AOI22X1_52 ( .A(_4426__bF_buf7), .B(_5179_), .C(_7998_), .D(_7931_), .Y(_81__5_) );
OAI21X1 OAI21X1_1378 ( .A(_7624__bF_buf2), .B(_10734__6_), .C(cpu_state_5_bF_buf1_), .Y(_7999_) );
OAI21X1 OAI21X1_1379 ( .A(_7629__bF_buf1), .B(_7631__bF_buf0), .C(_7999_), .Y(_8000_) );
INVX1 INVX1_658 ( .A(_7928_), .Y(_8001_) );
NAND2X1 NAND2X1_484 ( .A(_8001_), .B(_7924_), .Y(_8002_) );
OAI21X1 OAI21X1_1380 ( .A(_5179_), .B(_7926_), .C(_8002_), .Y(_8003_) );
NAND2X1 NAND2X1_485 ( .A(_10734__6_), .B(decoded_imm_6_), .Y(_8004_) );
INVX1 INVX1_659 ( .A(decoded_imm_6_), .Y(_8005_) );
NAND2X1 NAND2X1_486 ( .A(_5174_), .B(_8005_), .Y(_8006_) );
NAND2X1 NAND2X1_487 ( .A(_8004_), .B(_8006_), .Y(_8007_) );
XNOR2X1 XNOR2X1_5 ( .A(_8003_), .B(_8007_), .Y(_8008_) );
NOR2X1 NOR2X1_602 ( .A(_7624__bF_buf1), .B(_7999_), .Y(_8009_) );
OAI21X1 OAI21X1_1381 ( .A(_8008_), .B(_8009_), .C(_8000_), .Y(_8010_) );
NAND2X1 NAND2X1_488 ( .A(cpuregs_6_[6]), .B(decoded_rs1_1_bF_buf31_), .Y(_8011_) );
OAI21X1 OAI21X1_1382 ( .A(_5709_), .B(decoded_rs1_1_bF_buf30_), .C(_8011_), .Y(_8012_) );
MUX2X1 MUX2X1_150 ( .A(cpuregs_7_[6]), .B(cpuregs_5_[6]), .S(decoded_rs1_1_bF_buf29_), .Y(_8013_) );
OAI21X1 OAI21X1_1383 ( .A(_8013_), .B(_7569__bF_buf24), .C(decoded_rs1_2_bF_buf9_), .Y(_8014_) );
AOI21X1 AOI21X1_351 ( .A(_7569__bF_buf23), .B(_8012_), .C(_8014_), .Y(_8015_) );
MUX2X1 MUX2X1_151 ( .A(cpuregs_2_[6]), .B(cpuregs_0_[6]), .S(decoded_rs1_1_bF_buf28_), .Y(_8016_) );
NOR2X1 NOR2X1_603 ( .A(decoded_rs1_0_bF_buf16_), .B(_8016_), .Y(_8017_) );
MUX2X1 MUX2X1_152 ( .A(cpuregs_3_[6]), .B(cpuregs_1_[6]), .S(decoded_rs1_1_bF_buf27_), .Y(_8018_) );
OAI21X1 OAI21X1_1384 ( .A(_8018_), .B(_7569__bF_buf22), .C(_7560__bF_buf1), .Y(_8019_) );
OAI21X1 OAI21X1_1385 ( .A(_8019_), .B(_8017_), .C(_7552__bF_buf3), .Y(_8020_) );
NOR2X1 NOR2X1_604 ( .A(_8015_), .B(_8020_), .Y(_8021_) );
NAND2X1 NAND2X1_489 ( .A(cpuregs_22_[6]), .B(decoded_rs1_1_bF_buf26_), .Y(_8022_) );
OAI21X1 OAI21X1_1386 ( .A(_5978_), .B(decoded_rs1_1_bF_buf25_), .C(_8022_), .Y(_8023_) );
MUX2X1 MUX2X1_153 ( .A(cpuregs_23_[6]), .B(cpuregs_21_[6]), .S(decoded_rs1_1_bF_buf24_), .Y(_8024_) );
OAI21X1 OAI21X1_1387 ( .A(_8024_), .B(_7569__bF_buf21), .C(decoded_rs1_2_bF_buf8_), .Y(_8025_) );
AOI21X1 AOI21X1_352 ( .A(_7569__bF_buf20), .B(_8023_), .C(_8025_), .Y(_8026_) );
NAND2X1 NAND2X1_490 ( .A(_5970_), .B(_7569__bF_buf19), .Y(_8027_) );
OAI21X1 OAI21X1_1388 ( .A(cpuregs_17_[6]), .B(_7569__bF_buf18), .C(_8027_), .Y(_8028_) );
NAND2X1 NAND2X1_491 ( .A(_5973_), .B(_7569__bF_buf17), .Y(_8029_) );
OAI21X1 OAI21X1_1389 ( .A(cpuregs_19_[6]), .B(_7569__bF_buf16), .C(_8029_), .Y(_8030_) );
MUX2X1 MUX2X1_154 ( .A(_8030_), .B(_8028_), .S(decoded_rs1_1_bF_buf23_), .Y(_8031_) );
OAI21X1 OAI21X1_1390 ( .A(_8031_), .B(decoded_rs1_2_bF_buf7_), .C(decoded_rs1_4_bF_buf1_), .Y(_8032_) );
OAI21X1 OAI21X1_1391 ( .A(_8032_), .B(_8026_), .C(_7561__bF_buf2), .Y(_8033_) );
NOR2X1 NOR2X1_605 ( .A(_8021_), .B(_8033_), .Y(_8034_) );
OAI21X1 OAI21X1_1392 ( .A(_7560__bF_buf0), .B(cpuregs_14_[6]), .C(_7569__bF_buf15), .Y(_8035_) );
AOI21X1 AOI21X1_353 ( .A(_5942_), .B(_7560__bF_buf12), .C(_8035_), .Y(_8036_) );
NOR2X1 NOR2X1_606 ( .A(cpuregs_11_[6]), .B(decoded_rs1_2_bF_buf6_), .Y(_8037_) );
OAI21X1 OAI21X1_1393 ( .A(_7560__bF_buf11), .B(cpuregs_15_[6]), .C(decoded_rs1_0_bF_buf15_), .Y(_8038_) );
NOR2X1 NOR2X1_607 ( .A(_8037_), .B(_8038_), .Y(_8039_) );
OAI21X1 OAI21X1_1394 ( .A(_8036_), .B(_8039_), .C(decoded_rs1_1_bF_buf22_), .Y(_8040_) );
OAI21X1 OAI21X1_1395 ( .A(_7560__bF_buf10), .B(cpuregs_12_[6]), .C(_7569__bF_buf14), .Y(_8041_) );
AOI21X1 AOI21X1_354 ( .A(_4657_), .B(_7560__bF_buf9), .C(_8041_), .Y(_8042_) );
OAI21X1 OAI21X1_1396 ( .A(_7560__bF_buf8), .B(cpuregs_13_[6]), .C(decoded_rs1_0_bF_buf14_), .Y(_8043_) );
AOI21X1 AOI21X1_355 ( .A(_5939_), .B(_7560__bF_buf7), .C(_8043_), .Y(_8044_) );
OAI21X1 OAI21X1_1397 ( .A(_8042_), .B(_8044_), .C(_7556__bF_buf31), .Y(_8045_) );
AOI21X1 AOI21X1_356 ( .A(_8040_), .B(_8045_), .C(decoded_rs1_4_bF_buf0_), .Y(_8046_) );
AOI21X1 AOI21X1_357 ( .A(decoded_rs1_2_bF_buf5_), .B(_5965_), .C(decoded_rs1_0_bF_buf13_), .Y(_8047_) );
OAI21X1 OAI21X1_1398 ( .A(cpuregs_26_[6]), .B(decoded_rs1_2_bF_buf4_), .C(_8047_), .Y(_8048_) );
NOR2X1 NOR2X1_608 ( .A(cpuregs_27_[6]), .B(decoded_rs1_2_bF_buf3_), .Y(_8049_) );
OAI21X1 OAI21X1_1399 ( .A(_7560__bF_buf6), .B(cpuregs_31_[6]), .C(decoded_rs1_0_bF_buf12_), .Y(_8050_) );
OAI21X1 OAI21X1_1400 ( .A(_8049_), .B(_8050_), .C(_8048_), .Y(_8051_) );
AOI21X1 AOI21X1_358 ( .A(decoded_rs1_2_bF_buf2_), .B(_5962_), .C(decoded_rs1_0_bF_buf11_), .Y(_8052_) );
OAI21X1 OAI21X1_1401 ( .A(cpuregs_24_[6]), .B(decoded_rs1_2_bF_buf1_), .C(_8052_), .Y(_8053_) );
NOR2X1 NOR2X1_609 ( .A(cpuregs_25_[6]), .B(decoded_rs1_2_bF_buf0_), .Y(_8054_) );
OAI21X1 OAI21X1_1402 ( .A(_7560__bF_buf5), .B(cpuregs_29_[6]), .C(decoded_rs1_0_bF_buf10_), .Y(_8055_) );
OAI21X1 OAI21X1_1403 ( .A(_8054_), .B(_8055_), .C(_8053_), .Y(_8056_) );
MUX2X1 MUX2X1_155 ( .A(_8056_), .B(_8051_), .S(_7556__bF_buf30), .Y(_8057_) );
OAI21X1 OAI21X1_1404 ( .A(_8057_), .B(_7552__bF_buf2), .C(decoded_rs1_3_bF_buf1_), .Y(_8058_) );
OAI21X1 OAI21X1_1405 ( .A(_8058_), .B(_8046_), .C(_7587_), .Y(_8059_) );
OAI22X1 OAI22X1_129 ( .A(_4658_), .B(_7643_), .C(_8059_), .D(_8034_), .Y(_8060_) );
NOR2X1 NOR2X1_610 ( .A(_5179_), .B(_7700__bF_buf3), .Y(_8061_) );
NOR2X1 NOR2X1_611 ( .A(_8061_), .B(_4580__bF_buf1), .Y(_8062_) );
OAI21X1 OAI21X1_1406 ( .A(_7778_), .B(_7700__bF_buf2), .C(_10734__10_), .Y(_8063_) );
NOR2X1 NOR2X1_612 ( .A(_7841_), .B(_4579__bF_buf1), .Y(_8064_) );
AOI22X1 AOI22X1_53 ( .A(_8063_), .B(_8064_), .C(_8062_), .D(_7844_), .Y(_8065_) );
AOI21X1 AOI21X1_359 ( .A(_8065_), .B(_4584_), .C(_4426__bF_buf6), .Y(_8066_) );
AOI21X1 AOI21X1_360 ( .A(_7630_), .B(_7631__bF_buf5), .C(_7639_), .Y(_8067_) );
OAI21X1 OAI21X1_1407 ( .A(_8067_), .B(_5174_), .C(_8066_), .Y(_8068_) );
AOI21X1 AOI21X1_361 ( .A(cpu_state_2_bF_buf3_), .B(_8060_), .C(_8068_), .Y(_8069_) );
AOI22X1 AOI22X1_54 ( .A(_4426__bF_buf5), .B(_5174_), .C(_8010_), .D(_8069_), .Y(_81__6_) );
INVX1 INVX1_660 ( .A(decoded_imm_7_), .Y(_8070_) );
NOR2X1 NOR2X1_613 ( .A(_5173_), .B(_8070_), .Y(_8071_) );
NOR2X1 NOR2X1_614 ( .A(_10734__7_), .B(decoded_imm_7_), .Y(_8072_) );
NOR2X1 NOR2X1_615 ( .A(_8072_), .B(_8071_), .Y(_8073_) );
INVX1 INVX1_661 ( .A(_8007_), .Y(_8074_) );
NAND2X1 NAND2X1_492 ( .A(_8074_), .B(_8003_), .Y(_8075_) );
OAI21X1 OAI21X1_1408 ( .A(_5174_), .B(_8005_), .C(_8075_), .Y(_8076_) );
XOR2X1 XOR2X1_5 ( .A(_8076_), .B(_8073_), .Y(_8077_) );
AOI21X1 AOI21X1_362 ( .A(_5173_), .B(_7631__bF_buf4), .C(_7629__bF_buf0), .Y(_8078_) );
OAI21X1 OAI21X1_1409 ( .A(_8077_), .B(_7631__bF_buf3), .C(_8078_), .Y(_8079_) );
AOI21X1 AOI21X1_363 ( .A(_5173_), .B(_7623__bF_buf0), .C(_4587__bF_buf1), .Y(_8080_) );
OAI21X1 OAI21X1_1410 ( .A(_8077_), .B(_7623__bF_buf4), .C(_8080_), .Y(_8081_) );
INVX1 INVX1_662 ( .A(reg_pc_7_), .Y(_8082_) );
AND2X2 AND2X2_56 ( .A(cpuregs_17_[7]), .B(decoded_rs1_0_bF_buf9_), .Y(_8083_) );
OAI21X1 OAI21X1_1411 ( .A(_6015_), .B(decoded_rs1_0_bF_buf8_), .C(_7556__bF_buf29), .Y(_8084_) );
AOI21X1 AOI21X1_364 ( .A(cpuregs_19_[7]), .B(decoded_rs1_0_bF_buf7_), .C(_7556__bF_buf28), .Y(_8085_) );
OAI21X1 OAI21X1_1412 ( .A(_6018_), .B(decoded_rs1_0_bF_buf6_), .C(_8085_), .Y(_8086_) );
OAI21X1 OAI21X1_1413 ( .A(_8083_), .B(_8084_), .C(_8086_), .Y(_8087_) );
NAND2X1 NAND2X1_493 ( .A(_7560__bF_buf4), .B(_8087_), .Y(_8088_) );
NAND2X1 NAND2X1_494 ( .A(_6023_), .B(_7569__bF_buf13), .Y(_8089_) );
OAI21X1 OAI21X1_1414 ( .A(cpuregs_21_[7]), .B(_7569__bF_buf12), .C(_8089_), .Y(_8090_) );
NAND2X1 NAND2X1_495 ( .A(decoded_rs1_0_bF_buf5_), .B(_6026_), .Y(_8091_) );
OAI21X1 OAI21X1_1415 ( .A(cpuregs_22_[7]), .B(decoded_rs1_0_bF_buf4_), .C(_8091_), .Y(_8092_) );
MUX2X1 MUX2X1_156 ( .A(_8090_), .B(_8092_), .S(_7556__bF_buf27), .Y(_8093_) );
OAI21X1 OAI21X1_1416 ( .A(_7560__bF_buf3), .B(_8093_), .C(_8088_), .Y(_8094_) );
NOR2X1 NOR2X1_616 ( .A(_6032_), .B(_7569__bF_buf11), .Y(_8095_) );
INVX1 INVX1_663 ( .A(cpuregs_24_[7]), .Y(_8096_) );
OAI21X1 OAI21X1_1417 ( .A(_8096_), .B(decoded_rs1_0_bF_buf3_), .C(_7556__bF_buf26), .Y(_8097_) );
INVX1 INVX1_664 ( .A(cpuregs_26_[7]), .Y(_8098_) );
AOI21X1 AOI21X1_365 ( .A(cpuregs_27_[7]), .B(decoded_rs1_0_bF_buf2_), .C(_7556__bF_buf25), .Y(_8099_) );
OAI21X1 OAI21X1_1418 ( .A(_8098_), .B(decoded_rs1_0_bF_buf1_), .C(_8099_), .Y(_8100_) );
OAI21X1 OAI21X1_1419 ( .A(_8095_), .B(_8097_), .C(_8100_), .Y(_8101_) );
NAND2X1 NAND2X1_496 ( .A(_7560__bF_buf2), .B(_8101_), .Y(_8102_) );
NAND2X1 NAND2X1_497 ( .A(cpuregs_29_[7]), .B(decoded_rs1_0_bF_buf0_), .Y(_8103_) );
AOI21X1 AOI21X1_366 ( .A(cpuregs_28_[7]), .B(_7569__bF_buf10), .C(decoded_rs1_1_bF_buf21_), .Y(_8104_) );
NAND2X1 NAND2X1_498 ( .A(_6041_), .B(_7569__bF_buf9), .Y(_8105_) );
OAI21X1 OAI21X1_1420 ( .A(cpuregs_31_[7]), .B(_7569__bF_buf8), .C(_8105_), .Y(_8106_) );
AOI22X1 AOI22X1_55 ( .A(_8103_), .B(_8104_), .C(_8106_), .D(decoded_rs1_1_bF_buf20_), .Y(_8107_) );
OAI21X1 OAI21X1_1421 ( .A(_7560__bF_buf1), .B(_8107_), .C(_8102_), .Y(_8108_) );
MUX2X1 MUX2X1_157 ( .A(_8108_), .B(_8094_), .S(decoded_rs1_3_bF_buf0_), .Y(_8109_) );
OAI21X1 OAI21X1_1422 ( .A(_7560__bF_buf0), .B(cpuregs_13_[7]), .C(decoded_rs1_0_bF_buf57_), .Y(_8110_) );
AOI21X1 AOI21X1_367 ( .A(_5991_), .B(_7560__bF_buf12), .C(_8110_), .Y(_8111_) );
NOR2X1 NOR2X1_617 ( .A(cpuregs_8_[7]), .B(decoded_rs1_2_bF_buf12_), .Y(_8112_) );
OAI21X1 OAI21X1_1423 ( .A(_7560__bF_buf11), .B(cpuregs_12_[7]), .C(_7569__bF_buf7), .Y(_8113_) );
OAI21X1 OAI21X1_1424 ( .A(_8113_), .B(_8112_), .C(_7556__bF_buf24), .Y(_8114_) );
NOR2X1 NOR2X1_618 ( .A(cpuregs_11_[7]), .B(decoded_rs1_2_bF_buf11_), .Y(_8115_) );
OAI21X1 OAI21X1_1425 ( .A(_7560__bF_buf10), .B(cpuregs_15_[7]), .C(decoded_rs1_0_bF_buf56_), .Y(_8116_) );
NOR2X1 NOR2X1_619 ( .A(_8115_), .B(_8116_), .Y(_8117_) );
NOR2X1 NOR2X1_620 ( .A(cpuregs_10_[7]), .B(decoded_rs1_2_bF_buf10_), .Y(_8118_) );
OAI21X1 OAI21X1_1426 ( .A(_7560__bF_buf9), .B(cpuregs_14_[7]), .C(_7569__bF_buf6), .Y(_8119_) );
OAI21X1 OAI21X1_1427 ( .A(_8119_), .B(_8118_), .C(decoded_rs1_1_bF_buf19_), .Y(_8120_) );
OAI22X1 OAI22X1_130 ( .A(_8114_), .B(_8111_), .C(_8117_), .D(_8120_), .Y(_8121_) );
AND2X2 AND2X2_57 ( .A(_8121_), .B(decoded_rs1_3_bF_buf6_), .Y(_8122_) );
MUX2X1 MUX2X1_158 ( .A(cpuregs_2_[7]), .B(cpuregs_0_[7]), .S(decoded_rs1_1_bF_buf18_), .Y(_8123_) );
NOR2X1 NOR2X1_621 ( .A(decoded_rs1_0_bF_buf55_), .B(_8123_), .Y(_8124_) );
MUX2X1 MUX2X1_159 ( .A(cpuregs_3_[7]), .B(cpuregs_1_[7]), .S(decoded_rs1_1_bF_buf17_), .Y(_8125_) );
OAI21X1 OAI21X1_1428 ( .A(_8125_), .B(_7569__bF_buf5), .C(_7560__bF_buf8), .Y(_8126_) );
MUX2X1 MUX2X1_160 ( .A(cpuregs_6_[7]), .B(cpuregs_4_[7]), .S(decoded_rs1_1_bF_buf16_), .Y(_8127_) );
NOR2X1 NOR2X1_622 ( .A(decoded_rs1_0_bF_buf54_), .B(_8127_), .Y(_8128_) );
MUX2X1 MUX2X1_161 ( .A(cpuregs_7_[7]), .B(cpuregs_5_[7]), .S(decoded_rs1_1_bF_buf15_), .Y(_8129_) );
OAI21X1 OAI21X1_1429 ( .A(_8129_), .B(_7569__bF_buf4), .C(decoded_rs1_2_bF_buf9_), .Y(_8130_) );
OAI22X1 OAI22X1_131 ( .A(_8126_), .B(_8124_), .C(_8128_), .D(_8130_), .Y(_8131_) );
AND2X2 AND2X2_58 ( .A(_8131_), .B(_7561__bF_buf1), .Y(_8132_) );
OAI21X1 OAI21X1_1430 ( .A(_8122_), .B(_8132_), .C(_7552__bF_buf1), .Y(_8133_) );
OAI21X1 OAI21X1_1431 ( .A(_8109_), .B(_7552__bF_buf0), .C(_8133_), .Y(_8134_) );
OAI22X1 OAI22X1_132 ( .A(_8082_), .B(_7643_), .C(_8134_), .D(_7586__bF_buf2), .Y(_8135_) );
OAI21X1 OAI21X1_1432 ( .A(_7778_), .B(_7700__bF_buf1), .C(_10734__8_), .Y(_8136_) );
OAI21X1 OAI21X1_1433 ( .A(_7778_), .B(_7700__bF_buf0), .C(_10734__11_), .Y(_8137_) );
NOR2X1 NOR2X1_623 ( .A(_7908_), .B(_4579__bF_buf0), .Y(_8138_) );
INVX1 INVX1_665 ( .A(_7700__bF_buf5), .Y(_8139_) );
AOI21X1 AOI21X1_368 ( .A(_10734__6_), .B(_8139_), .C(_4580__bF_buf0), .Y(_8140_) );
AOI22X1 AOI22X1_56 ( .A(_8137_), .B(_8138_), .C(_8140_), .D(_8136_), .Y(_8141_) );
AOI21X1 AOI21X1_369 ( .A(_8141_), .B(_4584_), .C(_4426__bF_buf4), .Y(_8142_) );
OAI21X1 OAI21X1_1434 ( .A(_5173_), .B(_7640_), .C(_8142_), .Y(_8143_) );
AOI21X1 AOI21X1_370 ( .A(cpu_state_2_bF_buf2_), .B(_8135_), .C(_8143_), .Y(_8144_) );
AND2X2 AND2X2_59 ( .A(_8081_), .B(_8144_), .Y(_8145_) );
AOI22X1 AOI22X1_57 ( .A(_4426__bF_buf3), .B(_5173_), .C(_8145_), .D(_8079_), .Y(_81__7_) );
OAI21X1 OAI21X1_1435 ( .A(_7778_), .B(_7700__bF_buf4), .C(_10734__12_), .Y(_8146_) );
NOR2X1 NOR2X1_624 ( .A(_7992_), .B(_4579__bF_buf4), .Y(_8147_) );
AOI21X1 AOI21X1_371 ( .A(_10734__7_), .B(_8139_), .C(_4580__bF_buf4), .Y(_8148_) );
AOI22X1 AOI22X1_58 ( .A(_8146_), .B(_8147_), .C(_8148_), .D(_7990_), .Y(_8149_) );
AOI21X1 AOI21X1_372 ( .A(_8149_), .B(_4584_), .C(_4426__bF_buf2), .Y(_8150_) );
OAI21X1 OAI21X1_1436 ( .A(_7928_), .B(_7923_), .C(_7925_), .Y(_8151_) );
AND2X2 AND2X2_60 ( .A(_8074_), .B(_8073_), .Y(_8152_) );
INVX1 INVX1_666 ( .A(_8071_), .Y(_8153_) );
OAI21X1 OAI21X1_1437 ( .A(_8072_), .B(_8004_), .C(_8153_), .Y(_8154_) );
AOI21X1 AOI21X1_373 ( .A(_8151_), .B(_8152_), .C(_8154_), .Y(_8155_) );
NAND3X1 NAND3X1_34 ( .A(_7916_), .B(_8001_), .C(_8152_), .Y(_8156_) );
OAI21X1 OAI21X1_1438 ( .A(_8156_), .B(_7919_), .C(_8155_), .Y(_8157_) );
XOR2X1 XOR2X1_6 ( .A(_10734__8_), .B(decoded_imm_8_), .Y(_8158_) );
NOR2X1 NOR2X1_625 ( .A(_8158_), .B(_8157_), .Y(_8159_) );
NAND2X1 NAND2X1_499 ( .A(_8158_), .B(_8157_), .Y(_8160_) );
INVX1 INVX1_667 ( .A(_8160_), .Y(_8161_) );
OAI21X1 OAI21X1_1439 ( .A(_8161_), .B(_8159_), .C(_7632__bF_buf2), .Y(_8162_) );
AOI21X1 AOI21X1_374 ( .A(_5187_), .B(_7631__bF_buf2), .C(_7629__bF_buf3), .Y(_8163_) );
NAND2X1 NAND2X1_500 ( .A(_8163_), .B(_8162_), .Y(_8164_) );
OAI21X1 OAI21X1_1440 ( .A(_8161_), .B(_8159_), .C(_7624__bF_buf0), .Y(_8165_) );
AOI21X1 AOI21X1_375 ( .A(_5187_), .B(_7623__bF_buf3), .C(_4587__bF_buf0), .Y(_8166_) );
OAI21X1 OAI21X1_1441 ( .A(_6093_), .B(decoded_rs1_0_bF_buf53_), .C(_7556__bF_buf23), .Y(_8167_) );
AOI21X1 AOI21X1_376 ( .A(cpuregs_17_[8]), .B(decoded_rs1_0_bF_buf52_), .C(_8167_), .Y(_8168_) );
INVX1 INVX1_668 ( .A(cpuregs_19_[8]), .Y(_8169_) );
OAI21X1 OAI21X1_1442 ( .A(_8169_), .B(_7569__bF_buf3), .C(decoded_rs1_1_bF_buf14_), .Y(_8170_) );
AOI21X1 AOI21X1_377 ( .A(cpuregs_18_[8]), .B(_7569__bF_buf2), .C(_8170_), .Y(_8171_) );
OAI21X1 OAI21X1_1443 ( .A(_8168_), .B(_8171_), .C(_7560__bF_buf7), .Y(_8172_) );
OAI21X1 OAI21X1_1444 ( .A(_6101_), .B(decoded_rs1_0_bF_buf51_), .C(_7556__bF_buf22), .Y(_8173_) );
AOI21X1 AOI21X1_378 ( .A(cpuregs_21_[8]), .B(decoded_rs1_0_bF_buf50_), .C(_8173_), .Y(_8174_) );
OAI21X1 OAI21X1_1445 ( .A(_6104_), .B(_7569__bF_buf1), .C(decoded_rs1_1_bF_buf13_), .Y(_8175_) );
AOI21X1 AOI21X1_379 ( .A(cpuregs_22_[8]), .B(_7569__bF_buf0), .C(_8175_), .Y(_8176_) );
OAI21X1 OAI21X1_1446 ( .A(_8174_), .B(_8176_), .C(decoded_rs1_2_bF_buf8_), .Y(_8177_) );
AOI21X1 AOI21X1_380 ( .A(_8172_), .B(_8177_), .C(decoded_rs1_3_bF_buf5_), .Y(_8178_) );
AOI21X1 AOI21X1_381 ( .A(_6082_), .B(_7556__bF_buf21), .C(decoded_rs1_0_bF_buf49_), .Y(_8179_) );
OAI21X1 OAI21X1_1447 ( .A(cpuregs_26_[8]), .B(_7556__bF_buf20), .C(_8179_), .Y(_8180_) );
NOR2X1 NOR2X1_626 ( .A(cpuregs_27_[8]), .B(_7556__bF_buf19), .Y(_8181_) );
OAI21X1 OAI21X1_1448 ( .A(cpuregs_25_[8]), .B(decoded_rs1_1_bF_buf12_), .C(decoded_rs1_0_bF_buf48_), .Y(_8182_) );
OAI21X1 OAI21X1_1449 ( .A(_8181_), .B(_8182_), .C(_8180_), .Y(_8183_) );
AOI21X1 AOI21X1_382 ( .A(_6085_), .B(_7556__bF_buf18), .C(decoded_rs1_0_bF_buf47_), .Y(_8184_) );
OAI21X1 OAI21X1_1450 ( .A(cpuregs_30_[8]), .B(_7556__bF_buf17), .C(_8184_), .Y(_8185_) );
NOR2X1 NOR2X1_627 ( .A(cpuregs_31_[8]), .B(_7556__bF_buf16), .Y(_8186_) );
OAI21X1 OAI21X1_1451 ( .A(cpuregs_29_[8]), .B(decoded_rs1_1_bF_buf11_), .C(decoded_rs1_0_bF_buf46_), .Y(_8187_) );
OAI21X1 OAI21X1_1452 ( .A(_8186_), .B(_8187_), .C(_8185_), .Y(_8188_) );
MUX2X1 MUX2X1_162 ( .A(_8188_), .B(_8183_), .S(decoded_rs1_2_bF_buf7_), .Y(_8189_) );
AND2X2 AND2X2_61 ( .A(_8189_), .B(decoded_rs1_3_bF_buf4_), .Y(_8190_) );
OAI21X1 OAI21X1_1453 ( .A(_8190_), .B(_8178_), .C(decoded_rs1_4_bF_buf4_), .Y(_8191_) );
NOR2X1 NOR2X1_628 ( .A(cpuregs_1_[8]), .B(decoded_rs1_2_bF_buf6_), .Y(_8192_) );
OAI21X1 OAI21X1_1454 ( .A(_7560__bF_buf6), .B(cpuregs_5_[8]), .C(decoded_rs1_0_bF_buf45_), .Y(_8193_) );
NOR2X1 NOR2X1_629 ( .A(_8192_), .B(_8193_), .Y(_8194_) );
NOR2X1 NOR2X1_630 ( .A(cpuregs_0_[8]), .B(decoded_rs1_2_bF_buf5_), .Y(_8195_) );
OAI21X1 OAI21X1_1455 ( .A(_7560__bF_buf5), .B(cpuregs_4_[8]), .C(_7569__bF_buf48), .Y(_8196_) );
OAI21X1 OAI21X1_1456 ( .A(_8196_), .B(_8195_), .C(_7556__bF_buf15), .Y(_8197_) );
NOR2X1 NOR2X1_631 ( .A(cpuregs_3_[8]), .B(decoded_rs1_2_bF_buf4_), .Y(_8198_) );
OAI21X1 OAI21X1_1457 ( .A(_7560__bF_buf4), .B(cpuregs_7_[8]), .C(decoded_rs1_0_bF_buf44_), .Y(_8199_) );
NOR2X1 NOR2X1_632 ( .A(_8198_), .B(_8199_), .Y(_8200_) );
NOR2X1 NOR2X1_633 ( .A(cpuregs_2_[8]), .B(decoded_rs1_2_bF_buf3_), .Y(_8201_) );
OAI21X1 OAI21X1_1458 ( .A(_7560__bF_buf3), .B(cpuregs_6_[8]), .C(_7569__bF_buf47), .Y(_8202_) );
OAI21X1 OAI21X1_1459 ( .A(_8202_), .B(_8201_), .C(decoded_rs1_1_bF_buf10_), .Y(_8203_) );
OAI22X1 OAI22X1_133 ( .A(_8197_), .B(_8194_), .C(_8200_), .D(_8203_), .Y(_8204_) );
AND2X2 AND2X2_62 ( .A(_8204_), .B(_7561__bF_buf0), .Y(_8205_) );
NOR2X1 NOR2X1_634 ( .A(cpuregs_14_[8]), .B(_7556__bF_buf14), .Y(_8206_) );
OAI21X1 OAI21X1_1460 ( .A(cpuregs_12_[8]), .B(decoded_rs1_1_bF_buf9_), .C(_7569__bF_buf46), .Y(_8207_) );
NOR2X1 NOR2X1_635 ( .A(cpuregs_15_[8]), .B(_7556__bF_buf13), .Y(_8208_) );
OAI21X1 OAI21X1_1461 ( .A(cpuregs_13_[8]), .B(decoded_rs1_1_bF_buf8_), .C(decoded_rs1_0_bF_buf43_), .Y(_8209_) );
OAI22X1 OAI22X1_134 ( .A(_8206_), .B(_8207_), .C(_8208_), .D(_8209_), .Y(_8210_) );
AOI21X1 AOI21X1_383 ( .A(_4678_), .B(_7556__bF_buf12), .C(decoded_rs1_0_bF_buf42_), .Y(_8211_) );
OAI21X1 OAI21X1_1462 ( .A(cpuregs_10_[8]), .B(_7556__bF_buf11), .C(_8211_), .Y(_8212_) );
AOI21X1 AOI21X1_384 ( .A(_6070_), .B(_7556__bF_buf10), .C(_7569__bF_buf45), .Y(_8213_) );
OAI21X1 OAI21X1_1463 ( .A(cpuregs_11_[8]), .B(_7556__bF_buf9), .C(_8213_), .Y(_8214_) );
AND2X2 AND2X2_63 ( .A(_8212_), .B(_8214_), .Y(_8215_) );
OAI21X1 OAI21X1_1464 ( .A(_8215_), .B(decoded_rs1_2_bF_buf2_), .C(decoded_rs1_3_bF_buf3_), .Y(_8216_) );
AOI21X1 AOI21X1_385 ( .A(decoded_rs1_2_bF_buf1_), .B(_8210_), .C(_8216_), .Y(_8217_) );
OAI21X1 OAI21X1_1465 ( .A(_8217_), .B(_8205_), .C(_7552__bF_buf5), .Y(_8218_) );
NAND3X1 NAND3X1_35 ( .A(_7587_), .B(_8191_), .C(_8218_), .Y(_8219_) );
OAI21X1 OAI21X1_1466 ( .A(_4679_), .B(_7643_), .C(_8219_), .Y(_8220_) );
NAND2X1 NAND2X1_501 ( .A(cpu_state_2_bF_buf1_), .B(_8220_), .Y(_8221_) );
OAI21X1 OAI21X1_1467 ( .A(_5187_), .B(_7640_), .C(_8221_), .Y(_8222_) );
AOI21X1 AOI21X1_386 ( .A(_8165_), .B(_8166_), .C(_8222_), .Y(_8223_) );
AND2X2 AND2X2_64 ( .A(_8223_), .B(_8164_), .Y(_8224_) );
AOI22X1 AOI22X1_59 ( .A(_4426__bF_buf1), .B(_5187_), .C(_8224_), .D(_8150_), .Y(_81__8_) );
INVX1 INVX1_669 ( .A(decoded_imm_9_), .Y(_8225_) );
NOR2X1 NOR2X1_636 ( .A(_5107_), .B(_8225_), .Y(_8226_) );
NOR2X1 NOR2X1_637 ( .A(_10734__9_), .B(decoded_imm_9_), .Y(_8227_) );
NOR2X1 NOR2X1_638 ( .A(_8227_), .B(_8226_), .Y(_8228_) );
INVX1 INVX1_670 ( .A(_8228_), .Y(_8229_) );
INVX1 INVX1_671 ( .A(decoded_imm_8_), .Y(_8230_) );
OAI21X1 OAI21X1_1468 ( .A(_5187_), .B(_8230_), .C(_8160_), .Y(_8231_) );
XNOR2X1 XNOR2X1_6 ( .A(_8231_), .B(_8229_), .Y(_8232_) );
AOI21X1 AOI21X1_387 ( .A(_5107_), .B(_7631__bF_buf1), .C(_7629__bF_buf2), .Y(_8233_) );
OAI21X1 OAI21X1_1469 ( .A(_8232_), .B(_7631__bF_buf0), .C(_8233_), .Y(_8234_) );
AOI21X1 AOI21X1_388 ( .A(_5107_), .B(_7623__bF_buf2), .C(_4587__bF_buf3), .Y(_8235_) );
OAI21X1 OAI21X1_1470 ( .A(_8232_), .B(_7623__bF_buf1), .C(_8235_), .Y(_8236_) );
INVX1 INVX1_672 ( .A(reg_pc_9_), .Y(_8237_) );
OAI21X1 OAI21X1_1471 ( .A(_7560__bF_buf2), .B(cpuregs_13_[9]), .C(decoded_rs1_0_bF_buf41_), .Y(_8238_) );
AOI21X1 AOI21X1_389 ( .A(_6127_), .B(_7560__bF_buf1), .C(_8238_), .Y(_8239_) );
NOR2X1 NOR2X1_639 ( .A(cpuregs_8_[9]), .B(decoded_rs1_2_bF_buf0_), .Y(_8240_) );
OAI21X1 OAI21X1_1472 ( .A(_7560__bF_buf0), .B(cpuregs_12_[9]), .C(_7569__bF_buf44), .Y(_8241_) );
OAI21X1 OAI21X1_1473 ( .A(_8241_), .B(_8240_), .C(_7556__bF_buf8), .Y(_8242_) );
NOR2X1 NOR2X1_640 ( .A(cpuregs_11_[9]), .B(decoded_rs1_2_bF_buf12_), .Y(_8243_) );
OAI21X1 OAI21X1_1474 ( .A(_7560__bF_buf12), .B(cpuregs_15_[9]), .C(decoded_rs1_0_bF_buf40_), .Y(_8244_) );
NOR2X1 NOR2X1_641 ( .A(_8243_), .B(_8244_), .Y(_8245_) );
NOR2X1 NOR2X1_642 ( .A(cpuregs_10_[9]), .B(decoded_rs1_2_bF_buf11_), .Y(_8246_) );
OAI21X1 OAI21X1_1475 ( .A(_7560__bF_buf11), .B(cpuregs_14_[9]), .C(_7569__bF_buf43), .Y(_8247_) );
OAI21X1 OAI21X1_1476 ( .A(_8247_), .B(_8246_), .C(decoded_rs1_1_bF_buf7_), .Y(_8248_) );
OAI22X1 OAI22X1_135 ( .A(_8242_), .B(_8239_), .C(_8245_), .D(_8248_), .Y(_8249_) );
NAND2X1 NAND2X1_502 ( .A(decoded_rs1_3_bF_buf2_), .B(_8249_), .Y(_8250_) );
NAND2X1 NAND2X1_503 ( .A(_6113_), .B(_7569__bF_buf42), .Y(_8251_) );
OAI21X1 OAI21X1_1477 ( .A(cpuregs_1_[9]), .B(_7569__bF_buf41), .C(_8251_), .Y(_8252_) );
NAND2X1 NAND2X1_504 ( .A(_6116_), .B(_7569__bF_buf40), .Y(_8253_) );
OAI21X1 OAI21X1_1478 ( .A(cpuregs_3_[9]), .B(_7569__bF_buf39), .C(_8253_), .Y(_8254_) );
MUX2X1 MUX2X1_163 ( .A(_8254_), .B(_8252_), .S(decoded_rs1_1_bF_buf6_), .Y(_8255_) );
MUX2X1 MUX2X1_164 ( .A(cpuregs_6_[9]), .B(cpuregs_4_[9]), .S(decoded_rs1_1_bF_buf5_), .Y(_8256_) );
NOR2X1 NOR2X1_643 ( .A(decoded_rs1_0_bF_buf39_), .B(_8256_), .Y(_8257_) );
MUX2X1 MUX2X1_165 ( .A(cpuregs_7_[9]), .B(cpuregs_5_[9]), .S(decoded_rs1_1_bF_buf4_), .Y(_8258_) );
OAI21X1 OAI21X1_1479 ( .A(_8258_), .B(_7569__bF_buf38), .C(decoded_rs1_2_bF_buf10_), .Y(_8259_) );
OAI22X1 OAI22X1_136 ( .A(_8257_), .B(_8259_), .C(_8255_), .D(decoded_rs1_2_bF_buf9_), .Y(_8260_) );
NAND2X1 NAND2X1_505 ( .A(_7561__bF_buf6), .B(_8260_), .Y(_8261_) );
AOI21X1 AOI21X1_390 ( .A(_8250_), .B(_8261_), .C(decoded_rs1_4_bF_buf3_), .Y(_8262_) );
OAI21X1 OAI21X1_1480 ( .A(_7560__bF_buf10), .B(cpuregs_21_[9]), .C(decoded_rs1_0_bF_buf38_), .Y(_8263_) );
AOI21X1 AOI21X1_391 ( .A(_6157_), .B(_7560__bF_buf9), .C(_8263_), .Y(_8264_) );
NOR2X1 NOR2X1_644 ( .A(cpuregs_16_[9]), .B(decoded_rs1_2_bF_buf8_), .Y(_8265_) );
OAI21X1 OAI21X1_1481 ( .A(_7560__bF_buf8), .B(cpuregs_20_[9]), .C(_7569__bF_buf37), .Y(_8266_) );
OAI21X1 OAI21X1_1482 ( .A(_8266_), .B(_8265_), .C(_7556__bF_buf7), .Y(_8267_) );
OAI21X1 OAI21X1_1483 ( .A(_7560__bF_buf7), .B(cpuregs_23_[9]), .C(decoded_rs1_0_bF_buf37_), .Y(_8268_) );
AOI21X1 AOI21X1_392 ( .A(_6160_), .B(_7560__bF_buf6), .C(_8268_), .Y(_8269_) );
NOR2X1 NOR2X1_645 ( .A(cpuregs_18_[9]), .B(decoded_rs1_2_bF_buf7_), .Y(_8270_) );
OAI21X1 OAI21X1_1484 ( .A(_7560__bF_buf5), .B(cpuregs_22_[9]), .C(_7569__bF_buf36), .Y(_8271_) );
OAI21X1 OAI21X1_1485 ( .A(_8271_), .B(_8270_), .C(decoded_rs1_1_bF_buf3_), .Y(_8272_) );
OAI22X1 OAI22X1_137 ( .A(_8267_), .B(_8264_), .C(_8269_), .D(_8272_), .Y(_8273_) );
OAI21X1 OAI21X1_1486 ( .A(cpuregs_25_[9]), .B(decoded_rs1_1_bF_buf2_), .C(decoded_rs1_0_bF_buf36_), .Y(_8274_) );
AOI21X1 AOI21X1_393 ( .A(_6145_), .B(decoded_rs1_1_bF_buf1_), .C(_8274_), .Y(_8275_) );
NOR2X1 NOR2X1_646 ( .A(cpuregs_26_[9]), .B(_7556__bF_buf6), .Y(_8276_) );
OAI21X1 OAI21X1_1487 ( .A(cpuregs_24_[9]), .B(decoded_rs1_1_bF_buf0_), .C(_7569__bF_buf35), .Y(_8277_) );
OAI21X1 OAI21X1_1488 ( .A(_8276_), .B(_8277_), .C(_7560__bF_buf4), .Y(_8278_) );
OAI21X1 OAI21X1_1489 ( .A(cpuregs_29_[9]), .B(decoded_rs1_1_bF_buf44_), .C(decoded_rs1_0_bF_buf35_), .Y(_8279_) );
AOI21X1 AOI21X1_394 ( .A(_6152_), .B(decoded_rs1_1_bF_buf43_), .C(_8279_), .Y(_8280_) );
NOR2X1 NOR2X1_647 ( .A(cpuregs_30_[9]), .B(_7556__bF_buf5), .Y(_8281_) );
OAI21X1 OAI21X1_1490 ( .A(cpuregs_28_[9]), .B(decoded_rs1_1_bF_buf42_), .C(_7569__bF_buf34), .Y(_8282_) );
OAI21X1 OAI21X1_1491 ( .A(_8281_), .B(_8282_), .C(decoded_rs1_2_bF_buf6_), .Y(_8283_) );
OAI22X1 OAI22X1_138 ( .A(_8278_), .B(_8275_), .C(_8280_), .D(_8283_), .Y(_8284_) );
MUX2X1 MUX2X1_166 ( .A(_8273_), .B(_8284_), .S(_7561__bF_buf5), .Y(_8285_) );
OAI21X1 OAI21X1_1492 ( .A(_8285_), .B(_7552__bF_buf4), .C(_7587_), .Y(_8286_) );
OAI22X1 OAI22X1_139 ( .A(_8237_), .B(_7643_), .C(_8262_), .D(_8286_), .Y(_8287_) );
OAI21X1 OAI21X1_1493 ( .A(_7778_), .B(_7700__bF_buf3), .C(_10734__13_), .Y(_8288_) );
NOR2X1 NOR2X1_648 ( .A(_8061_), .B(_4579__bF_buf3), .Y(_8289_) );
NOR2X1 NOR2X1_649 ( .A(_5187_), .B(_7700__bF_buf2), .Y(_8290_) );
NOR2X1 NOR2X1_650 ( .A(_8290_), .B(_4580__bF_buf3), .Y(_8291_) );
AOI22X1 AOI22X1_60 ( .A(_8288_), .B(_8289_), .C(_8291_), .D(_8063_), .Y(_8292_) );
AOI21X1 AOI21X1_395 ( .A(_8292_), .B(_4584_), .C(_4426__bF_buf0), .Y(_8293_) );
OAI21X1 OAI21X1_1494 ( .A(_5107_), .B(_7640_), .C(_8293_), .Y(_8294_) );
AOI21X1 AOI21X1_396 ( .A(cpu_state_2_bF_buf0_), .B(_8287_), .C(_8294_), .Y(_8295_) );
AND2X2 AND2X2_65 ( .A(_8236_), .B(_8295_), .Y(_8296_) );
AOI22X1 AOI22X1_61 ( .A(_4426__bF_buf11), .B(_5107_), .C(_8296_), .D(_8234_), .Y(_81__9_) );
NAND2X1 NAND2X1_506 ( .A(_10734__8_), .B(decoded_imm_8_), .Y(_8297_) );
INVX1 INVX1_673 ( .A(_8226_), .Y(_8298_) );
OAI21X1 OAI21X1_1495 ( .A(_8227_), .B(_8297_), .C(_8298_), .Y(_8299_) );
INVX1 INVX1_674 ( .A(_8299_), .Y(_8300_) );
OAI21X1 OAI21X1_1496 ( .A(_8160_), .B(_8229_), .C(_8300_), .Y(_8301_) );
INVX1 INVX1_675 ( .A(_8301_), .Y(_8302_) );
NAND2X1 NAND2X1_507 ( .A(_10734__10_), .B(decoded_imm_10_), .Y(_8303_) );
INVX1 INVX1_676 ( .A(decoded_imm_10_), .Y(_8304_) );
NAND2X1 NAND2X1_508 ( .A(_5121_), .B(_8304_), .Y(_8305_) );
NAND2X1 NAND2X1_509 ( .A(_8303_), .B(_8305_), .Y(_8306_) );
OR2X2 OR2X2_6 ( .A(_8302_), .B(_8306_), .Y(_8307_) );
NAND2X1 NAND2X1_510 ( .A(_8306_), .B(_8302_), .Y(_8308_) );
AND2X2 AND2X2_66 ( .A(_8307_), .B(_8308_), .Y(_8309_) );
AOI21X1 AOI21X1_397 ( .A(_5121_), .B(_7631__bF_buf5), .C(_7629__bF_buf1), .Y(_8310_) );
OAI21X1 OAI21X1_1497 ( .A(_8309_), .B(_7631__bF_buf4), .C(_8310_), .Y(_8311_) );
INVX1 INVX1_677 ( .A(_8309_), .Y(_8312_) );
OAI21X1 OAI21X1_1498 ( .A(_7624__bF_buf4), .B(_10734__10_), .C(cpu_state_5_bF_buf0_), .Y(_8313_) );
AOI21X1 AOI21X1_398 ( .A(_7624__bF_buf3), .B(_8312_), .C(_8313_), .Y(_8314_) );
NOR2X1 NOR2X1_651 ( .A(cpuregs_1_[10]), .B(decoded_rs1_2_bF_buf5_), .Y(_8315_) );
OAI21X1 OAI21X1_1499 ( .A(_7560__bF_buf3), .B(cpuregs_5_[10]), .C(decoded_rs1_0_bF_buf34_), .Y(_8316_) );
NOR2X1 NOR2X1_652 ( .A(_8315_), .B(_8316_), .Y(_8317_) );
NOR2X1 NOR2X1_653 ( .A(cpuregs_0_[10]), .B(decoded_rs1_2_bF_buf4_), .Y(_8318_) );
OAI21X1 OAI21X1_1500 ( .A(_7560__bF_buf2), .B(cpuregs_4_[10]), .C(_7569__bF_buf33), .Y(_8319_) );
OAI21X1 OAI21X1_1501 ( .A(_8319_), .B(_8318_), .C(_7556__bF_buf4), .Y(_8320_) );
NOR2X1 NOR2X1_654 ( .A(cpuregs_3_[10]), .B(decoded_rs1_2_bF_buf3_), .Y(_8321_) );
OAI21X1 OAI21X1_1502 ( .A(_7560__bF_buf1), .B(cpuregs_7_[10]), .C(decoded_rs1_0_bF_buf33_), .Y(_8322_) );
NOR2X1 NOR2X1_655 ( .A(_8321_), .B(_8322_), .Y(_8323_) );
NOR2X1 NOR2X1_656 ( .A(cpuregs_2_[10]), .B(decoded_rs1_2_bF_buf2_), .Y(_8324_) );
OAI21X1 OAI21X1_1503 ( .A(_7560__bF_buf0), .B(cpuregs_6_[10]), .C(_7569__bF_buf32), .Y(_8325_) );
OAI21X1 OAI21X1_1504 ( .A(_8325_), .B(_8324_), .C(decoded_rs1_1_bF_buf41_), .Y(_8326_) );
OAI22X1 OAI22X1_140 ( .A(_8320_), .B(_8317_), .C(_8323_), .D(_8326_), .Y(_8327_) );
AND2X2 AND2X2_67 ( .A(_8327_), .B(_7561__bF_buf4), .Y(_8328_) );
NOR2X1 NOR2X1_657 ( .A(cpuregs_14_[10]), .B(_7556__bF_buf3), .Y(_8329_) );
OAI21X1 OAI21X1_1505 ( .A(cpuregs_12_[10]), .B(decoded_rs1_1_bF_buf40_), .C(_7569__bF_buf31), .Y(_8330_) );
NOR2X1 NOR2X1_658 ( .A(cpuregs_15_[10]), .B(_7556__bF_buf2), .Y(_8331_) );
OAI21X1 OAI21X1_1506 ( .A(cpuregs_13_[10]), .B(decoded_rs1_1_bF_buf39_), .C(decoded_rs1_0_bF_buf32_), .Y(_8332_) );
OAI22X1 OAI22X1_141 ( .A(_8329_), .B(_8330_), .C(_8331_), .D(_8332_), .Y(_8333_) );
AOI21X1 AOI21X1_399 ( .A(_4697_), .B(_7556__bF_buf1), .C(decoded_rs1_0_bF_buf31_), .Y(_8334_) );
OAI21X1 OAI21X1_1507 ( .A(cpuregs_10_[10]), .B(_7556__bF_buf0), .C(_8334_), .Y(_8335_) );
AOI21X1 AOI21X1_400 ( .A(_6177_), .B(_7556__bF_buf42), .C(_7569__bF_buf30), .Y(_8336_) );
OAI21X1 OAI21X1_1508 ( .A(cpuregs_11_[10]), .B(_7556__bF_buf41), .C(_8336_), .Y(_8337_) );
AND2X2 AND2X2_68 ( .A(_8335_), .B(_8337_), .Y(_8338_) );
OAI21X1 OAI21X1_1509 ( .A(_8338_), .B(decoded_rs1_2_bF_buf1_), .C(decoded_rs1_3_bF_buf1_), .Y(_8339_) );
AOI21X1 AOI21X1_401 ( .A(decoded_rs1_2_bF_buf0_), .B(_8333_), .C(_8339_), .Y(_8340_) );
OAI21X1 OAI21X1_1510 ( .A(_8340_), .B(_8328_), .C(_7552__bF_buf3), .Y(_8341_) );
INVX1 INVX1_678 ( .A(cpuregs_16_[10]), .Y(_8342_) );
OAI21X1 OAI21X1_1511 ( .A(_8342_), .B(decoded_rs1_0_bF_buf30_), .C(_7556__bF_buf40), .Y(_8343_) );
AOI21X1 AOI21X1_402 ( .A(cpuregs_17_[10]), .B(decoded_rs1_0_bF_buf29_), .C(_8343_), .Y(_8344_) );
INVX1 INVX1_679 ( .A(cpuregs_19_[10]), .Y(_8345_) );
OAI21X1 OAI21X1_1512 ( .A(_8345_), .B(_7569__bF_buf29), .C(decoded_rs1_1_bF_buf38_), .Y(_8346_) );
AOI21X1 AOI21X1_403 ( .A(cpuregs_18_[10]), .B(_7569__bF_buf28), .C(_8346_), .Y(_8347_) );
OAI21X1 OAI21X1_1513 ( .A(_8347_), .B(_8344_), .C(_7560__bF_buf12), .Y(_8348_) );
OAI21X1 OAI21X1_1514 ( .A(_6207_), .B(decoded_rs1_0_bF_buf28_), .C(_7556__bF_buf39), .Y(_8349_) );
AOI21X1 AOI21X1_404 ( .A(cpuregs_21_[10]), .B(decoded_rs1_0_bF_buf27_), .C(_8349_), .Y(_8350_) );
OAI21X1 OAI21X1_1515 ( .A(_6210_), .B(_7569__bF_buf27), .C(decoded_rs1_1_bF_buf37_), .Y(_8351_) );
AOI21X1 AOI21X1_405 ( .A(cpuregs_22_[10]), .B(_7569__bF_buf26), .C(_8351_), .Y(_8352_) );
OAI21X1 OAI21X1_1516 ( .A(_8352_), .B(_8350_), .C(decoded_rs1_2_bF_buf12_), .Y(_8353_) );
AND2X2 AND2X2_69 ( .A(_8348_), .B(_8353_), .Y(_8354_) );
AOI21X1 AOI21X1_406 ( .A(_6222_), .B(_7556__bF_buf38), .C(decoded_rs1_0_bF_buf26_), .Y(_8355_) );
OAI21X1 OAI21X1_1517 ( .A(cpuregs_30_[10]), .B(_7556__bF_buf37), .C(_8355_), .Y(_8356_) );
INVX1 INVX1_680 ( .A(cpuregs_29_[10]), .Y(_8357_) );
AOI21X1 AOI21X1_407 ( .A(_8357_), .B(_7556__bF_buf36), .C(_7569__bF_buf25), .Y(_8358_) );
OAI21X1 OAI21X1_1518 ( .A(cpuregs_31_[10]), .B(_7556__bF_buf35), .C(_8358_), .Y(_8359_) );
AOI21X1 AOI21X1_408 ( .A(_8356_), .B(_8359_), .C(_7560__bF_buf11), .Y(_8360_) );
OAI21X1 OAI21X1_1519 ( .A(cpuregs_24_[10]), .B(decoded_rs1_1_bF_buf36_), .C(_7569__bF_buf24), .Y(_8361_) );
AOI21X1 AOI21X1_409 ( .A(_6218_), .B(decoded_rs1_1_bF_buf35_), .C(_8361_), .Y(_8362_) );
INVX1 INVX1_681 ( .A(cpuregs_27_[10]), .Y(_8363_) );
OAI21X1 OAI21X1_1520 ( .A(cpuregs_25_[10]), .B(decoded_rs1_1_bF_buf34_), .C(decoded_rs1_0_bF_buf25_), .Y(_8364_) );
AOI21X1 AOI21X1_410 ( .A(_8363_), .B(decoded_rs1_1_bF_buf33_), .C(_8364_), .Y(_8365_) );
OAI21X1 OAI21X1_1521 ( .A(_8362_), .B(_8365_), .C(_7560__bF_buf10), .Y(_8366_) );
NAND2X1 NAND2X1_511 ( .A(decoded_rs1_3_bF_buf0_), .B(_8366_), .Y(_8367_) );
OAI22X1 OAI22X1_142 ( .A(_8360_), .B(_8367_), .C(_8354_), .D(decoded_rs1_3_bF_buf6_), .Y(_8368_) );
AOI21X1 AOI21X1_411 ( .A(decoded_rs1_4_bF_buf2_), .B(_8368_), .C(_7586__bF_buf1), .Y(_8369_) );
AOI22X1 AOI22X1_62 ( .A(reg_pc_10_), .B(_7551__bF_buf1), .C(_8369_), .D(_8341_), .Y(_8370_) );
INVX1 INVX1_682 ( .A(_8137_), .Y(_8371_) );
NOR2X1 NOR2X1_659 ( .A(_5203_), .B(_7698__bF_buf2), .Y(_8372_) );
OAI21X1 OAI21X1_1522 ( .A(_5174_), .B(_7700__bF_buf1), .C(_4580__bF_buf2), .Y(_8373_) );
OAI21X1 OAI21X1_1523 ( .A(_5107_), .B(_7700__bF_buf0), .C(_4579__bF_buf2), .Y(_8374_) );
OAI22X1 OAI22X1_143 ( .A(_8371_), .B(_8374_), .C(_8373_), .D(_8372_), .Y(_8375_) );
OAI21X1 OAI21X1_1524 ( .A(_7697__bF_buf2), .B(_8375_), .C(resetn_bF_buf11), .Y(_8376_) );
AOI21X1 AOI21X1_412 ( .A(_10734__10_), .B(_7639_), .C(_8376_), .Y(_8377_) );
OAI21X1 OAI21X1_1525 ( .A(_8370_), .B(_4538__bF_buf4), .C(_8377_), .Y(_8378_) );
NOR2X1 NOR2X1_660 ( .A(_8378_), .B(_8314_), .Y(_8379_) );
AOI22X1 AOI22X1_63 ( .A(_4426__bF_buf10), .B(_5121_), .C(_8379_), .D(_8311_), .Y(_81__10_) );
OAI21X1 OAI21X1_1526 ( .A(_8302_), .B(_8306_), .C(_8303_), .Y(_8380_) );
XNOR2X1 XNOR2X1_7 ( .A(_10734__11_), .B(decoded_imm_11_), .Y(_8381_) );
XNOR2X1 XNOR2X1_8 ( .A(_8380_), .B(_8381_), .Y(_8382_) );
AOI21X1 AOI21X1_413 ( .A(_5117_), .B(_7623__bF_buf0), .C(_4587__bF_buf2), .Y(_8383_) );
OAI21X1 OAI21X1_1527 ( .A(_8382_), .B(_7623__bF_buf4), .C(_8383_), .Y(_8384_) );
INVX1 INVX1_683 ( .A(_8382_), .Y(_8385_) );
OAI21X1 OAI21X1_1528 ( .A(_7632__bF_buf1), .B(_10734__11_), .C(_7630_), .Y(_8386_) );
AOI21X1 AOI21X1_414 ( .A(_7632__bF_buf0), .B(_8385_), .C(_8386_), .Y(_8387_) );
AND2X2 AND2X2_70 ( .A(cpuregs_17_[11]), .B(decoded_rs1_0_bF_buf24_), .Y(_8388_) );
OAI21X1 OAI21X1_1529 ( .A(_6279_), .B(decoded_rs1_0_bF_buf23_), .C(_7556__bF_buf34), .Y(_8389_) );
AND2X2 AND2X2_71 ( .A(_7569__bF_buf23), .B(cpuregs_18_[11]), .Y(_8390_) );
OAI21X1 OAI21X1_1530 ( .A(_6282_), .B(_7569__bF_buf22), .C(decoded_rs1_1_bF_buf32_), .Y(_8391_) );
OAI22X1 OAI22X1_144 ( .A(_8389_), .B(_8388_), .C(_8391_), .D(_8390_), .Y(_8392_) );
NOR2X1 NOR2X1_661 ( .A(decoded_rs1_2_bF_buf11_), .B(_8392_), .Y(_8393_) );
AND2X2 AND2X2_72 ( .A(cpuregs_21_[11]), .B(decoded_rs1_0_bF_buf22_), .Y(_8394_) );
OAI21X1 OAI21X1_1531 ( .A(_6287_), .B(decoded_rs1_0_bF_buf21_), .C(_7556__bF_buf33), .Y(_8395_) );
NOR2X1 NOR2X1_662 ( .A(decoded_rs1_0_bF_buf20_), .B(_6290_), .Y(_8396_) );
INVX1 INVX1_684 ( .A(cpuregs_23_[11]), .Y(_8397_) );
OAI21X1 OAI21X1_1532 ( .A(_8397_), .B(_7569__bF_buf21), .C(decoded_rs1_1_bF_buf31_), .Y(_8398_) );
OAI22X1 OAI22X1_145 ( .A(_8395_), .B(_8394_), .C(_8398_), .D(_8396_), .Y(_8399_) );
OAI21X1 OAI21X1_1533 ( .A(_8399_), .B(_7560__bF_buf9), .C(_7561__bF_buf3), .Y(_8400_) );
NOR2X1 NOR2X1_663 ( .A(_8393_), .B(_8400_), .Y(_8401_) );
AOI21X1 AOI21X1_415 ( .A(_6268_), .B(_7556__bF_buf32), .C(decoded_rs1_0_bF_buf19_), .Y(_8402_) );
OAI21X1 OAI21X1_1534 ( .A(cpuregs_26_[11]), .B(_7556__bF_buf31), .C(_8402_), .Y(_8403_) );
NOR2X1 NOR2X1_664 ( .A(cpuregs_27_[11]), .B(_7556__bF_buf30), .Y(_8404_) );
OAI21X1 OAI21X1_1535 ( .A(cpuregs_25_[11]), .B(decoded_rs1_1_bF_buf30_), .C(decoded_rs1_0_bF_buf18_), .Y(_8405_) );
OAI21X1 OAI21X1_1536 ( .A(_8404_), .B(_8405_), .C(_8403_), .Y(_8406_) );
OAI21X1 OAI21X1_1537 ( .A(cpuregs_28_[11]), .B(decoded_rs1_1_bF_buf29_), .C(_7569__bF_buf20), .Y(_8407_) );
AOI21X1 AOI21X1_416 ( .A(_6274_), .B(decoded_rs1_1_bF_buf28_), .C(_8407_), .Y(_8408_) );
INVX1 INVX1_685 ( .A(cpuregs_31_[11]), .Y(_8409_) );
OAI21X1 OAI21X1_1538 ( .A(cpuregs_29_[11]), .B(decoded_rs1_1_bF_buf27_), .C(decoded_rs1_0_bF_buf17_), .Y(_8410_) );
AOI21X1 AOI21X1_417 ( .A(_8409_), .B(decoded_rs1_1_bF_buf26_), .C(_8410_), .Y(_8411_) );
OAI21X1 OAI21X1_1539 ( .A(_8408_), .B(_8411_), .C(decoded_rs1_2_bF_buf10_), .Y(_8412_) );
NAND2X1 NAND2X1_512 ( .A(decoded_rs1_3_bF_buf5_), .B(_8412_), .Y(_8413_) );
AOI21X1 AOI21X1_418 ( .A(_7560__bF_buf8), .B(_8406_), .C(_8413_), .Y(_8414_) );
OAI21X1 OAI21X1_1540 ( .A(_8414_), .B(_8401_), .C(decoded_rs1_4_bF_buf1_), .Y(_8415_) );
AOI21X1 AOI21X1_419 ( .A(_4704_), .B(_7556__bF_buf29), .C(decoded_rs1_0_bF_buf16_), .Y(_8416_) );
OAI21X1 OAI21X1_1541 ( .A(cpuregs_10_[11]), .B(_7556__bF_buf28), .C(_8416_), .Y(_8417_) );
AOI21X1 AOI21X1_420 ( .A(_6256_), .B(_7556__bF_buf27), .C(_7569__bF_buf19), .Y(_8418_) );
OAI21X1 OAI21X1_1542 ( .A(cpuregs_11_[11]), .B(_7556__bF_buf26), .C(_8418_), .Y(_8419_) );
AOI21X1 AOI21X1_421 ( .A(_8417_), .B(_8419_), .C(decoded_rs1_2_bF_buf9_), .Y(_8420_) );
AND2X2 AND2X2_73 ( .A(cpuregs_1_[11]), .B(decoded_rs1_0_bF_buf15_), .Y(_8421_) );
INVX1 INVX1_686 ( .A(cpuregs_0_[11]), .Y(_8422_) );
OAI21X1 OAI21X1_1543 ( .A(_8422_), .B(decoded_rs1_0_bF_buf14_), .C(_7556__bF_buf25), .Y(_8423_) );
NOR2X1 NOR2X1_665 ( .A(decoded_rs1_0_bF_buf13_), .B(_6236_), .Y(_8424_) );
INVX1 INVX1_687 ( .A(cpuregs_3_[11]), .Y(_8425_) );
OAI21X1 OAI21X1_1544 ( .A(_8425_), .B(_7569__bF_buf18), .C(decoded_rs1_1_bF_buf25_), .Y(_8426_) );
OAI22X1 OAI22X1_146 ( .A(_8423_), .B(_8421_), .C(_8426_), .D(_8424_), .Y(_8427_) );
NOR2X1 NOR2X1_666 ( .A(decoded_rs1_2_bF_buf8_), .B(_8427_), .Y(_8428_) );
AND2X2 AND2X2_74 ( .A(cpuregs_5_[11]), .B(decoded_rs1_0_bF_buf12_), .Y(_8429_) );
OAI21X1 OAI21X1_1545 ( .A(_5714_), .B(decoded_rs1_0_bF_buf11_), .C(_7556__bF_buf24), .Y(_8430_) );
NOR2X1 NOR2X1_667 ( .A(decoded_rs1_0_bF_buf10_), .B(_5289_), .Y(_8431_) );
INVX1 INVX1_688 ( .A(cpuregs_7_[11]), .Y(_8432_) );
OAI21X1 OAI21X1_1546 ( .A(_8432_), .B(_7569__bF_buf17), .C(decoded_rs1_1_bF_buf24_), .Y(_8433_) );
OAI22X1 OAI22X1_147 ( .A(_8430_), .B(_8429_), .C(_8433_), .D(_8431_), .Y(_8434_) );
OAI21X1 OAI21X1_1547 ( .A(_8434_), .B(_7560__bF_buf7), .C(_7561__bF_buf2), .Y(_8435_) );
INVX1 INVX1_689 ( .A(cpuregs_12_[11]), .Y(_8436_) );
AOI21X1 AOI21X1_422 ( .A(_8436_), .B(_7556__bF_buf23), .C(decoded_rs1_0_bF_buf9_), .Y(_8437_) );
OAI21X1 OAI21X1_1548 ( .A(cpuregs_14_[11]), .B(_7556__bF_buf22), .C(_8437_), .Y(_8438_) );
AOI21X1 AOI21X1_423 ( .A(_6249_), .B(_7556__bF_buf21), .C(_7569__bF_buf16), .Y(_8439_) );
OAI21X1 OAI21X1_1549 ( .A(cpuregs_15_[11]), .B(_7556__bF_buf20), .C(_8439_), .Y(_8440_) );
AND2X2 AND2X2_75 ( .A(_8438_), .B(_8440_), .Y(_8441_) );
OAI21X1 OAI21X1_1550 ( .A(_8441_), .B(_7560__bF_buf6), .C(decoded_rs1_3_bF_buf4_), .Y(_8442_) );
OAI22X1 OAI22X1_148 ( .A(_8428_), .B(_8435_), .C(_8442_), .D(_8420_), .Y(_8443_) );
AOI21X1 AOI21X1_424 ( .A(_7552__bF_buf2), .B(_8443_), .C(_7586__bF_buf0), .Y(_8444_) );
AOI22X1 AOI22X1_64 ( .A(reg_pc_11_), .B(_7551__bF_buf0), .C(_8444_), .D(_8415_), .Y(_8445_) );
INVX1 INVX1_690 ( .A(_8146_), .Y(_8446_) );
OAI21X1 OAI21X1_1551 ( .A(_5121_), .B(_7700__bF_buf5), .C(_4579__bF_buf1), .Y(_8447_) );
NOR2X1 NOR2X1_668 ( .A(_5087_), .B(_7698__bF_buf1), .Y(_8448_) );
OAI21X1 OAI21X1_1552 ( .A(_5173_), .B(_7700__bF_buf4), .C(_4580__bF_buf1), .Y(_8449_) );
OAI22X1 OAI22X1_149 ( .A(_8446_), .B(_8447_), .C(_8449_), .D(_8448_), .Y(_8450_) );
OAI21X1 OAI21X1_1553 ( .A(_7697__bF_buf1), .B(_8450_), .C(resetn_bF_buf10), .Y(_8451_) );
AOI21X1 AOI21X1_425 ( .A(_10734__11_), .B(_7639_), .C(_8451_), .Y(_8452_) );
OAI21X1 OAI21X1_1554 ( .A(_8445_), .B(_4538__bF_buf3), .C(_8452_), .Y(_8453_) );
NOR2X1 NOR2X1_669 ( .A(_8453_), .B(_8387_), .Y(_8454_) );
AOI22X1 AOI22X1_65 ( .A(_4426__bF_buf9), .B(_5117_), .C(_8454_), .D(_8384_), .Y(_81__11_) );
NAND2X1 NAND2X1_513 ( .A(_8158_), .B(_8228_), .Y(_8455_) );
NOR2X1 NOR2X1_670 ( .A(_8381_), .B(_8306_), .Y(_8456_) );
INVX1 INVX1_691 ( .A(_8456_), .Y(_8457_) );
NOR2X1 NOR2X1_671 ( .A(_8455_), .B(_8457_), .Y(_8458_) );
INVX1 INVX1_692 ( .A(decoded_imm_11_), .Y(_8459_) );
OAI21X1 OAI21X1_1555 ( .A(_5117_), .B(_8459_), .C(_8303_), .Y(_8460_) );
OAI21X1 OAI21X1_1556 ( .A(_10734__11_), .B(decoded_imm_11_), .C(_8460_), .Y(_8461_) );
OAI21X1 OAI21X1_1557 ( .A(_8457_), .B(_8300_), .C(_8461_), .Y(_8462_) );
AOI21X1 AOI21X1_426 ( .A(_8458_), .B(_8157_), .C(_8462_), .Y(_8463_) );
NAND2X1 NAND2X1_514 ( .A(_10734__12_), .B(decoded_imm_12_), .Y(_8464_) );
INVX1 INVX1_693 ( .A(decoded_imm_12_), .Y(_8465_) );
NAND2X1 NAND2X1_515 ( .A(_5197_), .B(_8465_), .Y(_8466_) );
AND2X2 AND2X2_76 ( .A(_8466_), .B(_8464_), .Y(_8467_) );
INVX1 INVX1_694 ( .A(_8467_), .Y(_8468_) );
OR2X2 OR2X2_7 ( .A(_8463_), .B(_8468_), .Y(_8469_) );
NAND2X1 NAND2X1_516 ( .A(_8468_), .B(_8463_), .Y(_8470_) );
AND2X2 AND2X2_77 ( .A(_8469_), .B(_8470_), .Y(_8471_) );
AOI21X1 AOI21X1_427 ( .A(_5197_), .B(_7623__bF_buf3), .C(_4587__bF_buf1), .Y(_8472_) );
OAI21X1 OAI21X1_1558 ( .A(_8471_), .B(_7623__bF_buf2), .C(_8472_), .Y(_8473_) );
INVX1 INVX1_695 ( .A(_8471_), .Y(_8474_) );
OAI21X1 OAI21X1_1559 ( .A(_7632__bF_buf3), .B(_10734__12_), .C(_7630_), .Y(_8475_) );
AOI21X1 AOI21X1_428 ( .A(_7632__bF_buf2), .B(_8474_), .C(_8475_), .Y(_8476_) );
AND2X2 AND2X2_78 ( .A(cpuregs_1_[12]), .B(decoded_rs1_0_bF_buf8_), .Y(_8477_) );
INVX1 INVX1_696 ( .A(cpuregs_0_[12]), .Y(_8478_) );
OAI21X1 OAI21X1_1560 ( .A(_8478_), .B(decoded_rs1_0_bF_buf7_), .C(_7556__bF_buf19), .Y(_8479_) );
NOR2X1 NOR2X1_672 ( .A(decoded_rs1_0_bF_buf6_), .B(_6317_), .Y(_8480_) );
INVX1 INVX1_697 ( .A(cpuregs_3_[12]), .Y(_8481_) );
OAI21X1 OAI21X1_1561 ( .A(_8481_), .B(_7569__bF_buf15), .C(decoded_rs1_1_bF_buf23_), .Y(_8482_) );
OAI22X1 OAI22X1_150 ( .A(_8479_), .B(_8477_), .C(_8482_), .D(_8480_), .Y(_8483_) );
NOR2X1 NOR2X1_673 ( .A(decoded_rs1_2_bF_buf7_), .B(_8483_), .Y(_8484_) );
AND2X2 AND2X2_79 ( .A(cpuregs_5_[12]), .B(decoded_rs1_0_bF_buf5_), .Y(_8485_) );
INVX1 INVX1_698 ( .A(cpuregs_4_[12]), .Y(_8486_) );
OAI21X1 OAI21X1_1562 ( .A(_8486_), .B(decoded_rs1_0_bF_buf4_), .C(_7556__bF_buf18), .Y(_8487_) );
NOR2X1 NOR2X1_674 ( .A(decoded_rs1_0_bF_buf3_), .B(_6311_), .Y(_8488_) );
INVX1 INVX1_699 ( .A(cpuregs_7_[12]), .Y(_8489_) );
OAI21X1 OAI21X1_1563 ( .A(_8489_), .B(_7569__bF_buf14), .C(decoded_rs1_1_bF_buf22_), .Y(_8490_) );
OAI22X1 OAI22X1_151 ( .A(_8487_), .B(_8485_), .C(_8490_), .D(_8488_), .Y(_8491_) );
OAI21X1 OAI21X1_1564 ( .A(_8491_), .B(_7560__bF_buf5), .C(_7561__bF_buf1), .Y(_8492_) );
NOR2X1 NOR2X1_675 ( .A(_8484_), .B(_8492_), .Y(_8493_) );
NOR2X1 NOR2X1_676 ( .A(cpuregs_14_[12]), .B(_7556__bF_buf17), .Y(_8494_) );
OAI21X1 OAI21X1_1565 ( .A(cpuregs_12_[12]), .B(decoded_rs1_1_bF_buf21_), .C(_7569__bF_buf13), .Y(_8495_) );
NOR2X1 NOR2X1_677 ( .A(cpuregs_15_[12]), .B(_7556__bF_buf16), .Y(_8496_) );
OAI21X1 OAI21X1_1566 ( .A(cpuregs_13_[12]), .B(decoded_rs1_1_bF_buf20_), .C(decoded_rs1_0_bF_buf2_), .Y(_8497_) );
OAI22X1 OAI22X1_152 ( .A(_8494_), .B(_8495_), .C(_8496_), .D(_8497_), .Y(_8498_) );
NOR2X1 NOR2X1_678 ( .A(cpuregs_10_[12]), .B(_7556__bF_buf15), .Y(_8499_) );
OAI21X1 OAI21X1_1567 ( .A(cpuregs_8_[12]), .B(decoded_rs1_1_bF_buf19_), .C(_7569__bF_buf12), .Y(_8500_) );
NOR2X1 NOR2X1_679 ( .A(cpuregs_11_[12]), .B(_7556__bF_buf14), .Y(_8501_) );
OAI21X1 OAI21X1_1568 ( .A(cpuregs_9_[12]), .B(decoded_rs1_1_bF_buf18_), .C(decoded_rs1_0_bF_buf1_), .Y(_8502_) );
OAI22X1 OAI22X1_153 ( .A(_8499_), .B(_8500_), .C(_8501_), .D(_8502_), .Y(_8503_) );
MUX2X1 MUX2X1_167 ( .A(_8503_), .B(_8498_), .S(_7560__bF_buf4), .Y(_8504_) );
AND2X2 AND2X2_80 ( .A(_8504_), .B(decoded_rs1_3_bF_buf3_), .Y(_8505_) );
OAI21X1 OAI21X1_1569 ( .A(_8505_), .B(_8493_), .C(_7552__bF_buf1), .Y(_8506_) );
AND2X2 AND2X2_81 ( .A(cpuregs_29_[12]), .B(decoded_rs1_0_bF_buf0_), .Y(_8507_) );
OAI21X1 OAI21X1_1570 ( .A(_6347_), .B(decoded_rs1_0_bF_buf57_), .C(_7556__bF_buf13), .Y(_8508_) );
AND2X2 AND2X2_82 ( .A(_7569__bF_buf11), .B(cpuregs_30_[12]), .Y(_8509_) );
OAI21X1 OAI21X1_1571 ( .A(_6350_), .B(_7569__bF_buf10), .C(decoded_rs1_1_bF_buf17_), .Y(_8510_) );
OAI22X1 OAI22X1_154 ( .A(_8508_), .B(_8507_), .C(_8510_), .D(_8509_), .Y(_8511_) );
INVX1 INVX1_700 ( .A(cpuregs_26_[12]), .Y(_8512_) );
OAI21X1 OAI21X1_1572 ( .A(cpuregs_24_[12]), .B(decoded_rs1_1_bF_buf16_), .C(_7569__bF_buf9), .Y(_8513_) );
AOI21X1 AOI21X1_429 ( .A(_8512_), .B(decoded_rs1_1_bF_buf15_), .C(_8513_), .Y(_8514_) );
OAI21X1 OAI21X1_1573 ( .A(cpuregs_25_[12]), .B(decoded_rs1_1_bF_buf14_), .C(decoded_rs1_0_bF_buf56_), .Y(_8515_) );
AOI21X1 AOI21X1_430 ( .A(_6343_), .B(decoded_rs1_1_bF_buf13_), .C(_8515_), .Y(_8516_) );
OAI21X1 OAI21X1_1574 ( .A(_8514_), .B(_8516_), .C(_7560__bF_buf3), .Y(_8517_) );
OAI21X1 OAI21X1_1575 ( .A(_7560__bF_buf2), .B(_8511_), .C(_8517_), .Y(_8518_) );
AND2X2 AND2X2_83 ( .A(cpuregs_17_[12]), .B(decoded_rs1_0_bF_buf55_), .Y(_8519_) );
OAI21X1 OAI21X1_1576 ( .A(_6325_), .B(decoded_rs1_0_bF_buf54_), .C(_7556__bF_buf12), .Y(_8520_) );
AND2X2 AND2X2_84 ( .A(_7569__bF_buf8), .B(cpuregs_18_[12]), .Y(_8521_) );
OAI21X1 OAI21X1_1577 ( .A(_6328_), .B(_7569__bF_buf7), .C(decoded_rs1_1_bF_buf12_), .Y(_8522_) );
OAI22X1 OAI22X1_155 ( .A(_8520_), .B(_8519_), .C(_8522_), .D(_8521_), .Y(_8523_) );
NOR2X1 NOR2X1_680 ( .A(decoded_rs1_2_bF_buf6_), .B(_8523_), .Y(_8524_) );
AND2X2 AND2X2_85 ( .A(cpuregs_21_[12]), .B(decoded_rs1_0_bF_buf53_), .Y(_8525_) );
OAI21X1 OAI21X1_1578 ( .A(_6332_), .B(decoded_rs1_0_bF_buf52_), .C(_7556__bF_buf11), .Y(_8526_) );
NOR2X1 NOR2X1_681 ( .A(decoded_rs1_0_bF_buf51_), .B(_6335_), .Y(_8527_) );
INVX1 INVX1_701 ( .A(cpuregs_23_[12]), .Y(_8528_) );
OAI21X1 OAI21X1_1579 ( .A(_8528_), .B(_7569__bF_buf6), .C(decoded_rs1_1_bF_buf11_), .Y(_8529_) );
OAI22X1 OAI22X1_156 ( .A(_8526_), .B(_8525_), .C(_8529_), .D(_8527_), .Y(_8530_) );
OAI21X1 OAI21X1_1580 ( .A(_8530_), .B(_7560__bF_buf1), .C(_7561__bF_buf0), .Y(_8531_) );
OAI22X1 OAI22X1_157 ( .A(_8524_), .B(_8531_), .C(_8518_), .D(_7561__bF_buf6), .Y(_8532_) );
AOI21X1 AOI21X1_431 ( .A(decoded_rs1_4_bF_buf0_), .B(_8532_), .C(_7586__bF_buf3), .Y(_8533_) );
AOI22X1 AOI22X1_66 ( .A(reg_pc_12_), .B(_7551__bF_buf3), .C(_8533_), .D(_8506_), .Y(_8534_) );
INVX1 INVX1_702 ( .A(_8288_), .Y(_8535_) );
OAI21X1 OAI21X1_1581 ( .A(_5117_), .B(_7700__bF_buf3), .C(_4579__bF_buf0), .Y(_8536_) );
OAI21X1 OAI21X1_1582 ( .A(_7698__bF_buf0), .B(_5051_), .C(_4580__bF_buf0), .Y(_8537_) );
OAI22X1 OAI22X1_158 ( .A(_8535_), .B(_8536_), .C(_8537_), .D(_8290_), .Y(_8538_) );
OAI21X1 OAI21X1_1583 ( .A(_7697__bF_buf0), .B(_8538_), .C(resetn_bF_buf9), .Y(_8539_) );
AOI21X1 AOI21X1_432 ( .A(_10734__12_), .B(_7639_), .C(_8539_), .Y(_8540_) );
OAI21X1 OAI21X1_1584 ( .A(_8534_), .B(_4538__bF_buf2), .C(_8540_), .Y(_8541_) );
NOR2X1 NOR2X1_682 ( .A(_8541_), .B(_8476_), .Y(_8542_) );
AOI22X1 AOI22X1_67 ( .A(_4426__bF_buf8), .B(_5197_), .C(_8542_), .D(_8473_), .Y(_81__12_) );
INVX1 INVX1_703 ( .A(decoded_imm_13_), .Y(_8543_) );
NOR2X1 NOR2X1_683 ( .A(_5196_), .B(_8543_), .Y(_8544_) );
NOR2X1 NOR2X1_684 ( .A(_10734__13_), .B(decoded_imm_13_), .Y(_8545_) );
NOR2X1 NOR2X1_685 ( .A(_8545_), .B(_8544_), .Y(_8546_) );
OAI21X1 OAI21X1_1585 ( .A(_8463_), .B(_8468_), .C(_8464_), .Y(_8547_) );
NOR2X1 NOR2X1_686 ( .A(_8546_), .B(_8547_), .Y(_8548_) );
AND2X2 AND2X2_86 ( .A(_8547_), .B(_8546_), .Y(_8549_) );
OAI21X1 OAI21X1_1586 ( .A(_8549_), .B(_8548_), .C(_7632__bF_buf1), .Y(_8550_) );
AOI21X1 AOI21X1_433 ( .A(_5196_), .B(_7631__bF_buf3), .C(_7629__bF_buf0), .Y(_8551_) );
NAND2X1 NAND2X1_517 ( .A(_8551_), .B(_8550_), .Y(_8552_) );
OAI21X1 OAI21X1_1587 ( .A(_8549_), .B(_8548_), .C(_7624__bF_buf2), .Y(_8553_) );
AOI21X1 AOI21X1_434 ( .A(_5196_), .B(_7623__bF_buf1), .C(_4587__bF_buf0), .Y(_8554_) );
OAI21X1 OAI21X1_1588 ( .A(_6386_), .B(decoded_rs1_0_bF_buf50_), .C(_7556__bF_buf10), .Y(_8555_) );
AOI21X1 AOI21X1_435 ( .A(cpuregs_17_[13]), .B(decoded_rs1_0_bF_buf49_), .C(_8555_), .Y(_8556_) );
NAND2X1 NAND2X1_518 ( .A(_6389_), .B(_7569__bF_buf5), .Y(_8557_) );
OAI21X1 OAI21X1_1589 ( .A(cpuregs_19_[13]), .B(_7569__bF_buf4), .C(_8557_), .Y(_8558_) );
AOI21X1 AOI21X1_436 ( .A(decoded_rs1_1_bF_buf10_), .B(_8558_), .C(_8556_), .Y(_8559_) );
AND2X2 AND2X2_87 ( .A(cpuregs_21_[13]), .B(decoded_rs1_0_bF_buf48_), .Y(_8560_) );
OAI21X1 OAI21X1_1590 ( .A(_6394_), .B(decoded_rs1_0_bF_buf47_), .C(_7556__bF_buf9), .Y(_8561_) );
AOI21X1 AOI21X1_437 ( .A(cpuregs_23_[13]), .B(decoded_rs1_0_bF_buf46_), .C(_7556__bF_buf8), .Y(_8562_) );
OAI21X1 OAI21X1_1591 ( .A(_6397_), .B(decoded_rs1_0_bF_buf45_), .C(_8562_), .Y(_8563_) );
OAI21X1 OAI21X1_1592 ( .A(_8560_), .B(_8561_), .C(_8563_), .Y(_8564_) );
OAI21X1 OAI21X1_1593 ( .A(_8564_), .B(_7560__bF_buf0), .C(_7561__bF_buf5), .Y(_8565_) );
AOI21X1 AOI21X1_438 ( .A(_7560__bF_buf12), .B(_8559_), .C(_8565_), .Y(_8566_) );
NOR2X1 NOR2X1_687 ( .A(cpuregs_26_[13]), .B(_7556__bF_buf7), .Y(_8567_) );
OAI21X1 OAI21X1_1594 ( .A(cpuregs_24_[13]), .B(decoded_rs1_1_bF_buf9_), .C(_7569__bF_buf3), .Y(_8568_) );
NOR2X1 NOR2X1_688 ( .A(cpuregs_27_[13]), .B(_7556__bF_buf6), .Y(_8569_) );
OAI21X1 OAI21X1_1595 ( .A(cpuregs_25_[13]), .B(decoded_rs1_1_bF_buf8_), .C(decoded_rs1_0_bF_buf44_), .Y(_8570_) );
OAI22X1 OAI22X1_159 ( .A(_8567_), .B(_8568_), .C(_8569_), .D(_8570_), .Y(_8571_) );
INVX1 INVX1_704 ( .A(cpuregs_28_[13]), .Y(_8572_) );
AOI21X1 AOI21X1_439 ( .A(_8572_), .B(_7556__bF_buf5), .C(decoded_rs1_0_bF_buf43_), .Y(_8573_) );
OAI21X1 OAI21X1_1596 ( .A(cpuregs_30_[13]), .B(_7556__bF_buf4), .C(_8573_), .Y(_8574_) );
AOI21X1 AOI21X1_440 ( .A(_6409_), .B(_7556__bF_buf3), .C(_7569__bF_buf2), .Y(_8575_) );
OAI21X1 OAI21X1_1597 ( .A(cpuregs_31_[13]), .B(_7556__bF_buf2), .C(_8575_), .Y(_8576_) );
NAND3X1 NAND3X1_36 ( .A(decoded_rs1_2_bF_buf5_), .B(_8574_), .C(_8576_), .Y(_8577_) );
OAI21X1 OAI21X1_1598 ( .A(decoded_rs1_2_bF_buf4_), .B(_8571_), .C(_8577_), .Y(_8578_) );
AND2X2 AND2X2_88 ( .A(_8578_), .B(decoded_rs1_3_bF_buf2_), .Y(_8579_) );
OAI21X1 OAI21X1_1599 ( .A(_8579_), .B(_8566_), .C(decoded_rs1_4_bF_buf4_), .Y(_8580_) );
NOR2X1 NOR2X1_689 ( .A(cpuregs_1_[13]), .B(decoded_rs1_2_bF_buf3_), .Y(_8581_) );
OAI21X1 OAI21X1_1600 ( .A(_7560__bF_buf11), .B(cpuregs_5_[13]), .C(decoded_rs1_0_bF_buf42_), .Y(_8582_) );
NOR2X1 NOR2X1_690 ( .A(_8581_), .B(_8582_), .Y(_8583_) );
NOR2X1 NOR2X1_691 ( .A(cpuregs_0_[13]), .B(decoded_rs1_2_bF_buf2_), .Y(_8584_) );
OAI21X1 OAI21X1_1601 ( .A(_7560__bF_buf10), .B(cpuregs_4_[13]), .C(_7569__bF_buf1), .Y(_8585_) );
OAI21X1 OAI21X1_1602 ( .A(_8585_), .B(_8584_), .C(_7556__bF_buf1), .Y(_8586_) );
NOR2X1 NOR2X1_692 ( .A(_8583_), .B(_8586_), .Y(_8587_) );
INVX1 INVX1_705 ( .A(cpuregs_7_[13]), .Y(_8588_) );
AOI21X1 AOI21X1_441 ( .A(decoded_rs1_2_bF_buf1_), .B(_8588_), .C(_7569__bF_buf0), .Y(_8589_) );
OAI21X1 OAI21X1_1603 ( .A(cpuregs_3_[13]), .B(decoded_rs1_2_bF_buf0_), .C(_8589_), .Y(_8590_) );
OAI21X1 OAI21X1_1604 ( .A(_7560__bF_buf9), .B(cpuregs_6_[13]), .C(_7569__bF_buf48), .Y(_8591_) );
AOI21X1 AOI21X1_442 ( .A(_6378_), .B(_7560__bF_buf8), .C(_8591_), .Y(_8592_) );
NOR2X1 NOR2X1_693 ( .A(_7556__bF_buf0), .B(_8592_), .Y(_8593_) );
AOI21X1 AOI21X1_443 ( .A(_8590_), .B(_8593_), .C(_8587_), .Y(_8594_) );
INVX1 INVX1_706 ( .A(cpuregs_12_[13]), .Y(_8595_) );
AOI21X1 AOI21X1_444 ( .A(_8595_), .B(_7556__bF_buf42), .C(decoded_rs1_0_bF_buf41_), .Y(_8596_) );
OAI21X1 OAI21X1_1605 ( .A(cpuregs_14_[13]), .B(_7556__bF_buf41), .C(_8596_), .Y(_8597_) );
AOI21X1 AOI21X1_445 ( .A(_6366_), .B(_7556__bF_buf40), .C(_7569__bF_buf47), .Y(_8598_) );
OAI21X1 OAI21X1_1606 ( .A(cpuregs_15_[13]), .B(_7556__bF_buf39), .C(_8598_), .Y(_8599_) );
AOI21X1 AOI21X1_446 ( .A(_8597_), .B(_8599_), .C(_7560__bF_buf7), .Y(_8600_) );
AOI21X1 AOI21X1_447 ( .A(cpuregs_8_[13]), .B(_7569__bF_buf46), .C(decoded_rs1_1_bF_buf7_), .Y(_8601_) );
OAI21X1 OAI21X1_1607 ( .A(_6360_), .B(_7569__bF_buf45), .C(_8601_), .Y(_8602_) );
AND2X2 AND2X2_89 ( .A(_7569__bF_buf44), .B(cpuregs_10_[13]), .Y(_8603_) );
INVX1 INVX1_707 ( .A(cpuregs_11_[13]), .Y(_8604_) );
OAI21X1 OAI21X1_1608 ( .A(_8604_), .B(_7569__bF_buf43), .C(decoded_rs1_1_bF_buf6_), .Y(_8605_) );
OAI21X1 OAI21X1_1609 ( .A(_8603_), .B(_8605_), .C(_8602_), .Y(_8606_) );
OAI21X1 OAI21X1_1610 ( .A(_8606_), .B(decoded_rs1_2_bF_buf12_), .C(decoded_rs1_3_bF_buf1_), .Y(_8607_) );
OAI22X1 OAI22X1_160 ( .A(_8600_), .B(_8607_), .C(_8594_), .D(decoded_rs1_3_bF_buf0_), .Y(_8608_) );
AOI21X1 AOI21X1_448 ( .A(_7552__bF_buf0), .B(_8608_), .C(_7586__bF_buf2), .Y(_8609_) );
AOI22X1 AOI22X1_68 ( .A(reg_pc_13_), .B(_7551__bF_buf2), .C(_8609_), .D(_8580_), .Y(_8610_) );
NOR2X1 NOR2X1_694 ( .A(_5107_), .B(_7700__bF_buf2), .Y(_8611_) );
OAI21X1 OAI21X1_1611 ( .A(_7698__bF_buf4), .B(_5057_), .C(_4580__bF_buf4), .Y(_8612_) );
OAI21X1 OAI21X1_1612 ( .A(_5197_), .B(_7700__bF_buf1), .C(_4579__bF_buf4), .Y(_8613_) );
OAI22X1 OAI22X1_161 ( .A(_8372_), .B(_8613_), .C(_8612_), .D(_8611_), .Y(_8614_) );
OAI21X1 OAI21X1_1613 ( .A(_7697__bF_buf3), .B(_8614_), .C(resetn_bF_buf8), .Y(_8615_) );
AOI21X1 AOI21X1_449 ( .A(_10734__13_), .B(_7639_), .C(_8615_), .Y(_8616_) );
OAI21X1 OAI21X1_1614 ( .A(_8610_), .B(_4538__bF_buf1), .C(_8616_), .Y(_8617_) );
AOI21X1 AOI21X1_450 ( .A(_8554_), .B(_8553_), .C(_8617_), .Y(_8618_) );
AOI22X1 AOI22X1_69 ( .A(_4426__bF_buf7), .B(_5196_), .C(_8618_), .D(_8552_), .Y(_81__13_) );
NAND2X1 NAND2X1_519 ( .A(_8467_), .B(_8546_), .Y(_8619_) );
INVX1 INVX1_708 ( .A(_8464_), .Y(_8620_) );
AOI21X1 AOI21X1_451 ( .A(_8620_), .B(_8546_), .C(_8544_), .Y(_8621_) );
OAI21X1 OAI21X1_1615 ( .A(_8463_), .B(_8619_), .C(_8621_), .Y(_8622_) );
INVX1 INVX1_709 ( .A(decoded_imm_14_), .Y(_8623_) );
NOR2X1 NOR2X1_695 ( .A(_5203_), .B(_8623_), .Y(_8624_) );
NOR2X1 NOR2X1_696 ( .A(_10734__14_), .B(decoded_imm_14_), .Y(_8625_) );
NOR2X1 NOR2X1_697 ( .A(_8625_), .B(_8624_), .Y(_8626_) );
NOR2X1 NOR2X1_698 ( .A(_8626_), .B(_8622_), .Y(_8627_) );
AND2X2 AND2X2_90 ( .A(_8622_), .B(_8626_), .Y(_8628_) );
OAI21X1 OAI21X1_1616 ( .A(_8628_), .B(_8627_), .C(_7624__bF_buf1), .Y(_8629_) );
AOI21X1 AOI21X1_452 ( .A(_5203_), .B(_7623__bF_buf0), .C(_4587__bF_buf3), .Y(_8630_) );
NAND2X1 NAND2X1_520 ( .A(_8630_), .B(_8629_), .Y(_8631_) );
OAI21X1 OAI21X1_1617 ( .A(_8628_), .B(_8627_), .C(_7632__bF_buf0), .Y(_8632_) );
AOI21X1 AOI21X1_453 ( .A(_5203_), .B(_7631__bF_buf2), .C(_7629__bF_buf3), .Y(_8633_) );
INVX1 INVX1_710 ( .A(cpuregs_10_[14]), .Y(_8634_) );
OAI21X1 OAI21X1_1618 ( .A(_7560__bF_buf6), .B(cpuregs_14_[14]), .C(_7569__bF_buf42), .Y(_8635_) );
AOI21X1 AOI21X1_454 ( .A(_8634_), .B(_7560__bF_buf5), .C(_8635_), .Y(_8636_) );
INVX1 INVX1_711 ( .A(cpuregs_11_[14]), .Y(_8637_) );
OAI21X1 OAI21X1_1619 ( .A(_7560__bF_buf4), .B(cpuregs_15_[14]), .C(decoded_rs1_0_bF_buf40_), .Y(_8638_) );
AOI21X1 AOI21X1_455 ( .A(_8637_), .B(_7560__bF_buf3), .C(_8638_), .Y(_8639_) );
OAI21X1 OAI21X1_1620 ( .A(_8636_), .B(_8639_), .C(decoded_rs1_1_bF_buf5_), .Y(_8640_) );
NOR2X1 NOR2X1_699 ( .A(cpuregs_8_[14]), .B(decoded_rs1_2_bF_buf11_), .Y(_8641_) );
OAI21X1 OAI21X1_1621 ( .A(_7560__bF_buf2), .B(cpuregs_12_[14]), .C(_7569__bF_buf41), .Y(_8642_) );
NOR2X1 NOR2X1_700 ( .A(_8641_), .B(_8642_), .Y(_8643_) );
OAI21X1 OAI21X1_1622 ( .A(_7560__bF_buf1), .B(cpuregs_13_[14]), .C(decoded_rs1_0_bF_buf39_), .Y(_8644_) );
AOI21X1 AOI21X1_456 ( .A(_6468_), .B(_7560__bF_buf0), .C(_8644_), .Y(_8645_) );
OAI21X1 OAI21X1_1623 ( .A(_8645_), .B(_8643_), .C(_7556__bF_buf38), .Y(_8646_) );
NAND2X1 NAND2X1_521 ( .A(_8646_), .B(_8640_), .Y(_8647_) );
NOR2X1 NOR2X1_701 ( .A(_7561__bF_buf4), .B(_8647_), .Y(_8648_) );
INVX1 INVX1_712 ( .A(cpuregs_4_[14]), .Y(_8649_) );
OAI21X1 OAI21X1_1624 ( .A(_8649_), .B(decoded_rs1_0_bF_buf38_), .C(_7556__bF_buf37), .Y(_8650_) );
AOI21X1 AOI21X1_457 ( .A(cpuregs_5_[14]), .B(decoded_rs1_0_bF_buf37_), .C(_8650_), .Y(_8651_) );
INVX1 INVX1_713 ( .A(cpuregs_7_[14]), .Y(_8652_) );
OAI21X1 OAI21X1_1625 ( .A(_8652_), .B(_7569__bF_buf40), .C(decoded_rs1_1_bF_buf4_), .Y(_8653_) );
AOI21X1 AOI21X1_458 ( .A(cpuregs_6_[14]), .B(_7569__bF_buf39), .C(_8653_), .Y(_8654_) );
OAI21X1 OAI21X1_1626 ( .A(_8654_), .B(_8651_), .C(decoded_rs1_2_bF_buf10_), .Y(_8655_) );
INVX1 INVX1_714 ( .A(cpuregs_0_[14]), .Y(_8656_) );
OAI21X1 OAI21X1_1627 ( .A(_8656_), .B(decoded_rs1_0_bF_buf36_), .C(_7556__bF_buf36), .Y(_8657_) );
AOI21X1 AOI21X1_459 ( .A(cpuregs_1_[14]), .B(decoded_rs1_0_bF_buf35_), .C(_8657_), .Y(_8658_) );
INVX1 INVX1_715 ( .A(cpuregs_3_[14]), .Y(_8659_) );
OAI21X1 OAI21X1_1628 ( .A(_8659_), .B(_7569__bF_buf38), .C(decoded_rs1_1_bF_buf3_), .Y(_8660_) );
AOI21X1 AOI21X1_460 ( .A(cpuregs_2_[14]), .B(_7569__bF_buf37), .C(_8660_), .Y(_8661_) );
OAI21X1 OAI21X1_1629 ( .A(_8661_), .B(_8658_), .C(_7560__bF_buf12), .Y(_8662_) );
AOI21X1 AOI21X1_461 ( .A(_8655_), .B(_8662_), .C(decoded_rs1_3_bF_buf6_), .Y(_8663_) );
OAI21X1 OAI21X1_1630 ( .A(_8648_), .B(_8663_), .C(_7552__bF_buf5), .Y(_8664_) );
OAI21X1 OAI21X1_1631 ( .A(_6459_), .B(decoded_rs1_0_bF_buf34_), .C(_7556__bF_buf35), .Y(_8665_) );
AOI21X1 AOI21X1_462 ( .A(cpuregs_25_[14]), .B(decoded_rs1_0_bF_buf33_), .C(_8665_), .Y(_8666_) );
OAI21X1 OAI21X1_1632 ( .A(_6462_), .B(_7569__bF_buf36), .C(decoded_rs1_1_bF_buf2_), .Y(_8667_) );
AOI21X1 AOI21X1_463 ( .A(cpuregs_26_[14]), .B(_7569__bF_buf35), .C(_8667_), .Y(_8668_) );
OAI21X1 OAI21X1_1633 ( .A(_8668_), .B(_8666_), .C(_7560__bF_buf11), .Y(_8669_) );
OAI21X1 OAI21X1_1634 ( .A(_6451_), .B(decoded_rs1_0_bF_buf32_), .C(_7556__bF_buf34), .Y(_8670_) );
AOI21X1 AOI21X1_464 ( .A(cpuregs_29_[14]), .B(decoded_rs1_0_bF_buf31_), .C(_8670_), .Y(_8671_) );
OAI21X1 OAI21X1_1635 ( .A(_6454_), .B(_7569__bF_buf34), .C(decoded_rs1_1_bF_buf1_), .Y(_8672_) );
AOI21X1 AOI21X1_465 ( .A(cpuregs_30_[14]), .B(_7569__bF_buf33), .C(_8672_), .Y(_8673_) );
OAI21X1 OAI21X1_1636 ( .A(_8673_), .B(_8671_), .C(decoded_rs1_2_bF_buf9_), .Y(_8674_) );
AND2X2 AND2X2_91 ( .A(_8669_), .B(_8674_), .Y(_8675_) );
NOR2X1 NOR2X1_702 ( .A(_6426_), .B(_7569__bF_buf32), .Y(_8676_) );
OAI21X1 OAI21X1_1637 ( .A(_6423_), .B(decoded_rs1_0_bF_buf30_), .C(_7556__bF_buf33), .Y(_8677_) );
NOR2X1 NOR2X1_703 ( .A(decoded_rs1_0_bF_buf29_), .B(_6430_), .Y(_8678_) );
OAI21X1 OAI21X1_1638 ( .A(_6433_), .B(_7569__bF_buf31), .C(decoded_rs1_1_bF_buf0_), .Y(_8679_) );
OAI22X1 OAI22X1_162 ( .A(_8677_), .B(_8676_), .C(_8679_), .D(_8678_), .Y(_8680_) );
INVX1 INVX1_716 ( .A(cpuregs_16_[14]), .Y(_8681_) );
NAND2X1 NAND2X1_522 ( .A(cpuregs_18_[14]), .B(decoded_rs1_1_bF_buf44_), .Y(_8682_) );
OAI21X1 OAI21X1_1639 ( .A(_8681_), .B(decoded_rs1_1_bF_buf43_), .C(_8682_), .Y(_8683_) );
NAND2X1 NAND2X1_523 ( .A(_7569__bF_buf30), .B(_8683_), .Y(_8684_) );
INVX1 INVX1_717 ( .A(cpuregs_17_[14]), .Y(_8685_) );
NAND2X1 NAND2X1_524 ( .A(cpuregs_19_[14]), .B(decoded_rs1_1_bF_buf42_), .Y(_8686_) );
OAI21X1 OAI21X1_1640 ( .A(_8685_), .B(decoded_rs1_1_bF_buf41_), .C(_8686_), .Y(_8687_) );
AOI21X1 AOI21X1_466 ( .A(decoded_rs1_0_bF_buf28_), .B(_8687_), .C(decoded_rs1_2_bF_buf8_), .Y(_8688_) );
AOI22X1 AOI22X1_70 ( .A(_8684_), .B(_8688_), .C(_8680_), .D(decoded_rs1_2_bF_buf7_), .Y(_8689_) );
MUX2X1 MUX2X1_168 ( .A(_8675_), .B(_8689_), .S(decoded_rs1_3_bF_buf5_), .Y(_8690_) );
AOI21X1 AOI21X1_467 ( .A(decoded_rs1_4_bF_buf3_), .B(_8690_), .C(_7586__bF_buf1), .Y(_8691_) );
AOI22X1 AOI22X1_71 ( .A(reg_pc_14_), .B(_7551__bF_buf1), .C(_8691_), .D(_8664_), .Y(_8692_) );
OAI21X1 OAI21X1_1641 ( .A(_5196_), .B(_7700__bF_buf0), .C(_4579__bF_buf3), .Y(_8693_) );
NOR2X1 NOR2X1_704 ( .A(_5045_), .B(_7698__bF_buf3), .Y(_8694_) );
OAI21X1 OAI21X1_1642 ( .A(_5121_), .B(_7700__bF_buf5), .C(_4580__bF_buf3), .Y(_8695_) );
OAI22X1 OAI22X1_163 ( .A(_8448_), .B(_8693_), .C(_8695_), .D(_8694_), .Y(_8696_) );
OAI21X1 OAI21X1_1643 ( .A(_7697__bF_buf2), .B(_8696_), .C(resetn_bF_buf7), .Y(_8697_) );
AOI21X1 AOI21X1_468 ( .A(_10734__14_), .B(_7639_), .C(_8697_), .Y(_8698_) );
OAI21X1 OAI21X1_1644 ( .A(_4538__bF_buf0), .B(_8692_), .C(_8698_), .Y(_8699_) );
AOI21X1 AOI21X1_469 ( .A(_8633_), .B(_8632_), .C(_8699_), .Y(_8700_) );
AOI22X1 AOI22X1_72 ( .A(_4426__bF_buf6), .B(_5203_), .C(_8700_), .D(_8631_), .Y(_81__14_) );
NOR2X1 NOR2X1_705 ( .A(_8624_), .B(_8628_), .Y(_8701_) );
XOR2X1 XOR2X1_7 ( .A(_10734__15_), .B(decoded_imm_15_), .Y(_8702_) );
XNOR2X1 XNOR2X1_9 ( .A(_8701_), .B(_8702_), .Y(_8703_) );
AOI21X1 AOI21X1_470 ( .A(_5087_), .B(_7623__bF_buf4), .C(_4587__bF_buf2), .Y(_8704_) );
OAI21X1 OAI21X1_1645 ( .A(_8703_), .B(_7623__bF_buf3), .C(_8704_), .Y(_8705_) );
AOI21X1 AOI21X1_471 ( .A(_5087_), .B(_7631__bF_buf1), .C(_7629__bF_buf2), .Y(_8706_) );
OAI21X1 OAI21X1_1646 ( .A(_8703_), .B(_7631__bF_buf0), .C(_8706_), .Y(_8707_) );
OAI21X1 OAI21X1_1647 ( .A(_6519_), .B(decoded_rs1_0_bF_buf27_), .C(_7556__bF_buf32), .Y(_8708_) );
AOI21X1 AOI21X1_472 ( .A(cpuregs_25_[15]), .B(decoded_rs1_0_bF_buf26_), .C(_8708_), .Y(_8709_) );
OAI21X1 OAI21X1_1648 ( .A(_6522_), .B(_7569__bF_buf29), .C(decoded_rs1_1_bF_buf40_), .Y(_8710_) );
AOI21X1 AOI21X1_473 ( .A(cpuregs_26_[15]), .B(_7569__bF_buf28), .C(_8710_), .Y(_8711_) );
OAI21X1 OAI21X1_1649 ( .A(_8709_), .B(_8711_), .C(_7560__bF_buf10), .Y(_8712_) );
OAI21X1 OAI21X1_1650 ( .A(_6511_), .B(decoded_rs1_0_bF_buf25_), .C(_7556__bF_buf31), .Y(_8713_) );
AOI21X1 AOI21X1_474 ( .A(cpuregs_29_[15]), .B(decoded_rs1_0_bF_buf24_), .C(_8713_), .Y(_8714_) );
OAI21X1 OAI21X1_1651 ( .A(_6514_), .B(_7569__bF_buf27), .C(decoded_rs1_1_bF_buf39_), .Y(_8715_) );
AOI21X1 AOI21X1_475 ( .A(cpuregs_30_[15]), .B(_7569__bF_buf26), .C(_8715_), .Y(_8716_) );
OAI21X1 OAI21X1_1652 ( .A(_8714_), .B(_8716_), .C(decoded_rs1_2_bF_buf6_), .Y(_8717_) );
AOI21X1 AOI21X1_476 ( .A(_8712_), .B(_8717_), .C(_7561__bF_buf3), .Y(_8718_) );
MUX2X1 MUX2X1_169 ( .A(cpuregs_22_[15]), .B(cpuregs_20_[15]), .S(decoded_rs1_1_bF_buf38_), .Y(_8719_) );
NAND2X1 NAND2X1_525 ( .A(cpuregs_23_[15]), .B(decoded_rs1_1_bF_buf37_), .Y(_8720_) );
OAI21X1 OAI21X1_1653 ( .A(_6534_), .B(decoded_rs1_1_bF_buf36_), .C(_8720_), .Y(_8721_) );
AOI21X1 AOI21X1_477 ( .A(decoded_rs1_0_bF_buf23_), .B(_8721_), .C(_7560__bF_buf9), .Y(_8722_) );
OAI21X1 OAI21X1_1654 ( .A(decoded_rs1_0_bF_buf22_), .B(_8719_), .C(_8722_), .Y(_8723_) );
MUX2X1 MUX2X1_170 ( .A(cpuregs_18_[15]), .B(cpuregs_16_[15]), .S(decoded_rs1_1_bF_buf35_), .Y(_8724_) );
NAND2X1 NAND2X1_526 ( .A(cpuregs_19_[15]), .B(decoded_rs1_1_bF_buf34_), .Y(_8725_) );
OAI21X1 OAI21X1_1655 ( .A(_6528_), .B(decoded_rs1_1_bF_buf33_), .C(_8725_), .Y(_8726_) );
AOI21X1 AOI21X1_478 ( .A(decoded_rs1_0_bF_buf21_), .B(_8726_), .C(decoded_rs1_2_bF_buf5_), .Y(_8727_) );
OAI21X1 OAI21X1_1656 ( .A(decoded_rs1_0_bF_buf20_), .B(_8724_), .C(_8727_), .Y(_8728_) );
AOI21X1 AOI21X1_479 ( .A(_8723_), .B(_8728_), .C(decoded_rs1_3_bF_buf4_), .Y(_8729_) );
OAI21X1 OAI21X1_1657 ( .A(_8718_), .B(_8729_), .C(decoded_rs1_4_bF_buf2_), .Y(_8730_) );
AOI21X1 AOI21X1_480 ( .A(_6503_), .B(_7556__bF_buf30), .C(_7569__bF_buf25), .Y(_8731_) );
OAI21X1 OAI21X1_1658 ( .A(cpuregs_15_[15]), .B(_7556__bF_buf29), .C(_8731_), .Y(_8732_) );
INVX1 INVX1_718 ( .A(cpuregs_12_[15]), .Y(_8733_) );
AOI21X1 AOI21X1_481 ( .A(_8733_), .B(_7556__bF_buf28), .C(decoded_rs1_0_bF_buf19_), .Y(_8734_) );
OAI21X1 OAI21X1_1659 ( .A(cpuregs_14_[15]), .B(_7556__bF_buf27), .C(_8734_), .Y(_8735_) );
NAND3X1 NAND3X1_37 ( .A(decoded_rs1_2_bF_buf4_), .B(_8732_), .C(_8735_), .Y(_8736_) );
NOR2X1 NOR2X1_706 ( .A(_6497_), .B(_7569__bF_buf24), .Y(_8737_) );
INVX1 INVX1_719 ( .A(cpuregs_8_[15]), .Y(_8738_) );
OAI21X1 OAI21X1_1660 ( .A(_8738_), .B(decoded_rs1_0_bF_buf18_), .C(_7556__bF_buf26), .Y(_8739_) );
INVX1 INVX1_720 ( .A(cpuregs_10_[15]), .Y(_8740_) );
AOI21X1 AOI21X1_482 ( .A(cpuregs_11_[15]), .B(decoded_rs1_0_bF_buf17_), .C(_7556__bF_buf25), .Y(_8741_) );
OAI21X1 OAI21X1_1661 ( .A(_8740_), .B(decoded_rs1_0_bF_buf16_), .C(_8741_), .Y(_8742_) );
OAI21X1 OAI21X1_1662 ( .A(_8737_), .B(_8739_), .C(_8742_), .Y(_8743_) );
AOI21X1 AOI21X1_483 ( .A(_7560__bF_buf8), .B(_8743_), .C(_7561__bF_buf2), .Y(_8744_) );
INVX1 INVX1_721 ( .A(cpuregs_7_[15]), .Y(_8745_) );
AOI21X1 AOI21X1_484 ( .A(decoded_rs1_2_bF_buf3_), .B(_8745_), .C(_7569__bF_buf23), .Y(_8746_) );
OAI21X1 OAI21X1_1663 ( .A(cpuregs_3_[15]), .B(decoded_rs1_2_bF_buf2_), .C(_8746_), .Y(_8747_) );
OAI21X1 OAI21X1_1664 ( .A(_7560__bF_buf7), .B(cpuregs_6_[15]), .C(_7569__bF_buf22), .Y(_8748_) );
AOI21X1 AOI21X1_485 ( .A(_6490_), .B(_7560__bF_buf6), .C(_8748_), .Y(_8749_) );
NOR2X1 NOR2X1_707 ( .A(_7556__bF_buf24), .B(_8749_), .Y(_8750_) );
NOR2X1 NOR2X1_708 ( .A(cpuregs_1_[15]), .B(decoded_rs1_2_bF_buf1_), .Y(_8751_) );
OAI21X1 OAI21X1_1665 ( .A(_7560__bF_buf5), .B(cpuregs_5_[15]), .C(decoded_rs1_0_bF_buf15_), .Y(_8752_) );
NOR2X1 NOR2X1_709 ( .A(_8751_), .B(_8752_), .Y(_8753_) );
NOR2X1 NOR2X1_710 ( .A(cpuregs_0_[15]), .B(decoded_rs1_2_bF_buf0_), .Y(_8754_) );
OAI21X1 OAI21X1_1666 ( .A(_7560__bF_buf4), .B(cpuregs_4_[15]), .C(_7569__bF_buf21), .Y(_8755_) );
OAI21X1 OAI21X1_1667 ( .A(_8755_), .B(_8754_), .C(_7556__bF_buf23), .Y(_8756_) );
OAI21X1 OAI21X1_1668 ( .A(_8756_), .B(_8753_), .C(_7561__bF_buf1), .Y(_8757_) );
AOI21X1 AOI21X1_486 ( .A(_8747_), .B(_8750_), .C(_8757_), .Y(_8758_) );
AOI21X1 AOI21X1_487 ( .A(_8736_), .B(_8744_), .C(_8758_), .Y(_8759_) );
AOI21X1 AOI21X1_488 ( .A(_7552__bF_buf4), .B(_8759_), .C(_7586__bF_buf0), .Y(_8760_) );
AOI22X1 AOI22X1_73 ( .A(reg_pc_15_), .B(_7551__bF_buf0), .C(_8760_), .D(_8730_), .Y(_8761_) );
NOR2X1 NOR2X1_711 ( .A(_4538__bF_buf4), .B(_8761_), .Y(_8762_) );
NOR2X1 NOR2X1_712 ( .A(_5117_), .B(_7700__bF_buf4), .Y(_8763_) );
OAI21X1 OAI21X1_1669 ( .A(instr_slli), .B(instr_sll), .C(_10734__14_), .Y(_8764_) );
OAI21X1 OAI21X1_1670 ( .A(_7698__bF_buf2), .B(_5051_), .C(_8764_), .Y(_8765_) );
OAI21X1 OAI21X1_1671 ( .A(_7698__bF_buf1), .B(_5040_), .C(_4580__bF_buf2), .Y(_8766_) );
OAI22X1 OAI22X1_164 ( .A(_4580__bF_buf1), .B(_8765_), .C(_8766_), .D(_8763_), .Y(_8767_) );
OAI21X1 OAI21X1_1672 ( .A(_7627_), .B(_5087_), .C(resetn_bF_buf6), .Y(_8768_) );
AOI21X1 AOI21X1_489 ( .A(_10734__15_), .B(_4597__bF_buf2), .C(_8768_), .Y(_8769_) );
OAI21X1 OAI21X1_1673 ( .A(_7697__bF_buf1), .B(_8767_), .C(_8769_), .Y(_8770_) );
NOR2X1 NOR2X1_713 ( .A(_8770_), .B(_8762_), .Y(_8771_) );
AND2X2 AND2X2_92 ( .A(_8707_), .B(_8771_), .Y(_8772_) );
AOI22X1 AOI22X1_74 ( .A(_4426__bF_buf5), .B(_5087_), .C(_8772_), .D(_8705_), .Y(_81__15_) );
NAND2X1 NAND2X1_527 ( .A(_8702_), .B(_8626_), .Y(_8773_) );
NOR2X1 NOR2X1_714 ( .A(_8773_), .B(_8619_), .Y(_8774_) );
INVX1 INVX1_722 ( .A(decoded_imm_15_), .Y(_8775_) );
NOR2X1 NOR2X1_715 ( .A(_5087_), .B(_8775_), .Y(_8776_) );
AOI21X1 AOI21X1_490 ( .A(_8624_), .B(_8702_), .C(_8776_), .Y(_8777_) );
OAI21X1 OAI21X1_1674 ( .A(_8621_), .B(_8773_), .C(_8777_), .Y(_8778_) );
AOI21X1 AOI21X1_491 ( .A(_8462_), .B(_8774_), .C(_8778_), .Y(_8779_) );
NAND3X1 NAND3X1_38 ( .A(_8458_), .B(_8774_), .C(_8157_), .Y(_8780_) );
AND2X2 AND2X2_93 ( .A(_8780_), .B(_8779_), .Y(_8781_) );
INVX1 INVX1_723 ( .A(decoded_imm_16_), .Y(_8782_) );
NOR2X1 NOR2X1_716 ( .A(_5051_), .B(_8782_), .Y(_8783_) );
INVX1 INVX1_724 ( .A(_8783_), .Y(_8784_) );
NAND2X1 NAND2X1_528 ( .A(_5051_), .B(_8782_), .Y(_8785_) );
NAND2X1 NAND2X1_529 ( .A(_8785_), .B(_8784_), .Y(_8786_) );
NOR2X1 NOR2X1_717 ( .A(_8786_), .B(_8781_), .Y(_8787_) );
INVX1 INVX1_725 ( .A(_8787_), .Y(_8788_) );
NAND2X1 NAND2X1_530 ( .A(_8786_), .B(_8781_), .Y(_8789_) );
AND2X2 AND2X2_94 ( .A(_8788_), .B(_8789_), .Y(_8790_) );
AOI21X1 AOI21X1_492 ( .A(_5051_), .B(_7631__bF_buf5), .C(_7629__bF_buf1), .Y(_8791_) );
OAI21X1 OAI21X1_1675 ( .A(_8790_), .B(_7631__bF_buf4), .C(_8791_), .Y(_8792_) );
INVX1 INVX1_726 ( .A(_8790_), .Y(_8793_) );
OAI21X1 OAI21X1_1676 ( .A(_7624__bF_buf0), .B(_10734__16_), .C(cpu_state_5_bF_buf3_), .Y(_8794_) );
AOI21X1 AOI21X1_493 ( .A(_7624__bF_buf4), .B(_8793_), .C(_8794_), .Y(_8795_) );
OAI21X1 OAI21X1_1677 ( .A(_6583_), .B(decoded_rs1_0_bF_buf14_), .C(_7556__bF_buf22), .Y(_8796_) );
AOI21X1 AOI21X1_494 ( .A(cpuregs_25_[16]), .B(decoded_rs1_0_bF_buf13_), .C(_8796_), .Y(_8797_) );
OAI21X1 OAI21X1_1678 ( .A(_6586_), .B(_7569__bF_buf20), .C(decoded_rs1_1_bF_buf32_), .Y(_8798_) );
AOI21X1 AOI21X1_495 ( .A(cpuregs_26_[16]), .B(_7569__bF_buf19), .C(_8798_), .Y(_8799_) );
OAI21X1 OAI21X1_1679 ( .A(_8799_), .B(_8797_), .C(_7560__bF_buf3), .Y(_8800_) );
INVX1 INVX1_727 ( .A(cpuregs_28_[16]), .Y(_8801_) );
OAI21X1 OAI21X1_1680 ( .A(_8801_), .B(decoded_rs1_0_bF_buf12_), .C(_7556__bF_buf21), .Y(_8802_) );
AOI21X1 AOI21X1_496 ( .A(cpuregs_29_[16]), .B(decoded_rs1_0_bF_buf11_), .C(_8802_), .Y(_8803_) );
OAI21X1 OAI21X1_1681 ( .A(_6578_), .B(_7569__bF_buf18), .C(decoded_rs1_1_bF_buf31_), .Y(_8804_) );
AOI21X1 AOI21X1_497 ( .A(cpuregs_30_[16]), .B(_7569__bF_buf17), .C(_8804_), .Y(_8805_) );
OAI21X1 OAI21X1_1682 ( .A(_8805_), .B(_8803_), .C(decoded_rs1_2_bF_buf12_), .Y(_8806_) );
AND2X2 AND2X2_95 ( .A(_8800_), .B(_8806_), .Y(_8807_) );
INVX1 INVX1_728 ( .A(cpuregs_11_[16]), .Y(_8808_) );
OAI21X1 OAI21X1_1683 ( .A(cpuregs_9_[16]), .B(decoded_rs1_1_bF_buf30_), .C(decoded_rs1_0_bF_buf10_), .Y(_8809_) );
AOI21X1 AOI21X1_498 ( .A(_8808_), .B(decoded_rs1_1_bF_buf29_), .C(_8809_), .Y(_8810_) );
NOR2X1 NOR2X1_718 ( .A(cpuregs_10_[16]), .B(_7556__bF_buf20), .Y(_8811_) );
OAI21X1 OAI21X1_1684 ( .A(cpuregs_8_[16]), .B(decoded_rs1_1_bF_buf28_), .C(_7569__bF_buf16), .Y(_8812_) );
OAI21X1 OAI21X1_1685 ( .A(_8811_), .B(_8812_), .C(_7560__bF_buf2), .Y(_8813_) );
INVX1 INVX1_729 ( .A(cpuregs_15_[16]), .Y(_8814_) );
OAI21X1 OAI21X1_1686 ( .A(cpuregs_13_[16]), .B(decoded_rs1_1_bF_buf27_), .C(decoded_rs1_0_bF_buf9_), .Y(_8815_) );
AOI21X1 AOI21X1_499 ( .A(_8814_), .B(decoded_rs1_1_bF_buf26_), .C(_8815_), .Y(_8816_) );
NOR2X1 NOR2X1_719 ( .A(cpuregs_14_[16]), .B(_7556__bF_buf19), .Y(_8817_) );
OAI21X1 OAI21X1_1687 ( .A(cpuregs_12_[16]), .B(decoded_rs1_1_bF_buf25_), .C(_7569__bF_buf15), .Y(_8818_) );
OAI21X1 OAI21X1_1688 ( .A(_8817_), .B(_8818_), .C(decoded_rs1_2_bF_buf11_), .Y(_8819_) );
OAI22X1 OAI22X1_165 ( .A(_8813_), .B(_8810_), .C(_8816_), .D(_8819_), .Y(_8820_) );
NAND2X1 NAND2X1_531 ( .A(_7552__bF_buf3), .B(_8820_), .Y(_8821_) );
OAI21X1 OAI21X1_1689 ( .A(_8807_), .B(_7552__bF_buf2), .C(_8821_), .Y(_8822_) );
NAND2X1 NAND2X1_532 ( .A(decoded_rs1_3_bF_buf3_), .B(_8822_), .Y(_8823_) );
INVX1 INVX1_730 ( .A(cpuregs_16_[16]), .Y(_8824_) );
NAND2X1 NAND2X1_533 ( .A(cpuregs_18_[16]), .B(decoded_rs1_1_bF_buf24_), .Y(_8825_) );
OAI21X1 OAI21X1_1690 ( .A(_8824_), .B(decoded_rs1_1_bF_buf23_), .C(_8825_), .Y(_8826_) );
NAND2X1 NAND2X1_534 ( .A(_7569__bF_buf14), .B(_8826_), .Y(_8827_) );
INVX1 INVX1_731 ( .A(cpuregs_17_[16]), .Y(_8828_) );
NAND2X1 NAND2X1_535 ( .A(cpuregs_19_[16]), .B(decoded_rs1_1_bF_buf22_), .Y(_8829_) );
OAI21X1 OAI21X1_1691 ( .A(_8828_), .B(decoded_rs1_1_bF_buf21_), .C(_8829_), .Y(_8830_) );
AOI21X1 AOI21X1_500 ( .A(decoded_rs1_0_bF_buf8_), .B(_8830_), .C(decoded_rs1_2_bF_buf10_), .Y(_8831_) );
NOR2X1 NOR2X1_720 ( .A(_6550_), .B(_7569__bF_buf13), .Y(_8832_) );
OAI21X1 OAI21X1_1692 ( .A(_6547_), .B(decoded_rs1_0_bF_buf7_), .C(_7556__bF_buf18), .Y(_8833_) );
NOR2X1 NOR2X1_721 ( .A(decoded_rs1_0_bF_buf6_), .B(_6554_), .Y(_8834_) );
OAI21X1 OAI21X1_1693 ( .A(_6557_), .B(_7569__bF_buf12), .C(decoded_rs1_1_bF_buf20_), .Y(_8835_) );
OAI22X1 OAI22X1_166 ( .A(_8833_), .B(_8832_), .C(_8835_), .D(_8834_), .Y(_8836_) );
AOI22X1 AOI22X1_75 ( .A(_8827_), .B(_8831_), .C(_8836_), .D(decoded_rs1_2_bF_buf9_), .Y(_8837_) );
NOR2X1 NOR2X1_722 ( .A(cpuregs_1_[16]), .B(decoded_rs1_2_bF_buf8_), .Y(_8838_) );
OAI21X1 OAI21X1_1694 ( .A(_7560__bF_buf1), .B(cpuregs_5_[16]), .C(decoded_rs1_0_bF_buf5_), .Y(_8839_) );
NOR2X1 NOR2X1_723 ( .A(_8838_), .B(_8839_), .Y(_8840_) );
NOR2X1 NOR2X1_724 ( .A(cpuregs_0_[16]), .B(decoded_rs1_2_bF_buf7_), .Y(_8841_) );
OAI21X1 OAI21X1_1695 ( .A(_7560__bF_buf0), .B(cpuregs_4_[16]), .C(_7569__bF_buf11), .Y(_8842_) );
OAI21X1 OAI21X1_1696 ( .A(_8842_), .B(_8841_), .C(_7556__bF_buf17), .Y(_8843_) );
NOR2X1 NOR2X1_725 ( .A(cpuregs_3_[16]), .B(decoded_rs1_2_bF_buf6_), .Y(_8844_) );
OAI21X1 OAI21X1_1697 ( .A(_7560__bF_buf12), .B(cpuregs_7_[16]), .C(decoded_rs1_0_bF_buf4_), .Y(_8845_) );
NOR2X1 NOR2X1_726 ( .A(_8844_), .B(_8845_), .Y(_8846_) );
NOR2X1 NOR2X1_727 ( .A(cpuregs_2_[16]), .B(decoded_rs1_2_bF_buf5_), .Y(_8847_) );
OAI21X1 OAI21X1_1698 ( .A(_7560__bF_buf11), .B(cpuregs_6_[16]), .C(_7569__bF_buf10), .Y(_8848_) );
OAI21X1 OAI21X1_1699 ( .A(_8848_), .B(_8847_), .C(decoded_rs1_1_bF_buf19_), .Y(_8849_) );
OAI22X1 OAI22X1_167 ( .A(_8843_), .B(_8840_), .C(_8846_), .D(_8849_), .Y(_8850_) );
NAND2X1 NAND2X1_536 ( .A(_7552__bF_buf1), .B(_8850_), .Y(_8851_) );
OAI21X1 OAI21X1_1700 ( .A(_7552__bF_buf0), .B(_8837_), .C(_8851_), .Y(_8852_) );
AOI21X1 AOI21X1_501 ( .A(_7561__bF_buf0), .B(_8852_), .C(_7586__bF_buf3), .Y(_8853_) );
AOI22X1 AOI22X1_76 ( .A(reg_pc_16_), .B(_7551__bF_buf3), .C(_8823_), .D(_8853_), .Y(_8854_) );
INVX1 INVX1_732 ( .A(_7627_), .Y(_8855_) );
OAI21X1 OAI21X1_1701 ( .A(_4597__bF_buf1), .B(_8855_), .C(_10734__16_), .Y(_8856_) );
OAI21X1 OAI21X1_1702 ( .A(_8854_), .B(_4538__bF_buf3), .C(_8856_), .Y(_8857_) );
NOR2X1 NOR2X1_728 ( .A(_8857_), .B(_8795_), .Y(_8858_) );
AND2X2 AND2X2_96 ( .A(_8858_), .B(_8792_), .Y(_8859_) );
OAI21X1 OAI21X1_1703 ( .A(instr_slli), .B(instr_sll), .C(_10734__15_), .Y(_8860_) );
OAI21X1 OAI21X1_1704 ( .A(_7698__bF_buf0), .B(_5057_), .C(_8860_), .Y(_8861_) );
NAND2X1 NAND2X1_537 ( .A(_4579__bF_buf2), .B(_8861_), .Y(_8862_) );
NOR2X1 NOR2X1_729 ( .A(_5197_), .B(_7700__bF_buf3), .Y(_8863_) );
NOR2X1 NOR2X1_730 ( .A(_5218_), .B(_7698__bF_buf4), .Y(_8864_) );
OAI21X1 OAI21X1_1705 ( .A(_8864_), .B(_8863_), .C(_4580__bF_buf0), .Y(_8865_) );
NAND2X1 NAND2X1_538 ( .A(_8862_), .B(_8865_), .Y(_8866_) );
AOI21X1 AOI21X1_502 ( .A(_8866_), .B(_4584_), .C(_4426__bF_buf4), .Y(_8867_) );
AOI22X1 AOI22X1_77 ( .A(_4426__bF_buf3), .B(_5051_), .C(_8859_), .D(_8867_), .Y(_81__16_) );
INVX1 INVX1_733 ( .A(decoded_imm_17_), .Y(_8868_) );
NOR2X1 NOR2X1_731 ( .A(_5057_), .B(_8868_), .Y(_8869_) );
NOR2X1 NOR2X1_732 ( .A(_10734__17_), .B(decoded_imm_17_), .Y(_8870_) );
OAI21X1 OAI21X1_1706 ( .A(_8869_), .B(_8870_), .C(_8784_), .Y(_8871_) );
NOR2X1 NOR2X1_733 ( .A(_8871_), .B(_8787_), .Y(_8872_) );
NOR2X1 NOR2X1_734 ( .A(_8870_), .B(_8869_), .Y(_8873_) );
NAND2X1 NAND2X1_539 ( .A(_8783_), .B(_8873_), .Y(_8874_) );
NAND3X1 NAND3X1_39 ( .A(_8784_), .B(_8785_), .C(_8873_), .Y(_8875_) );
OAI21X1 OAI21X1_1707 ( .A(_8781_), .B(_8875_), .C(_8874_), .Y(_8876_) );
OR2X2 OR2X2_8 ( .A(_8872_), .B(_8876_), .Y(_8877_) );
INVX1 INVX1_734 ( .A(_8877_), .Y(_8878_) );
AOI21X1 AOI21X1_503 ( .A(_5057_), .B(_7631__bF_buf3), .C(_7629__bF_buf0), .Y(_8879_) );
OAI21X1 OAI21X1_1708 ( .A(_8878_), .B(_7631__bF_buf2), .C(_8879_), .Y(_8880_) );
OAI21X1 OAI21X1_1709 ( .A(_7624__bF_buf3), .B(_10734__17_), .C(cpu_state_5_bF_buf2_), .Y(_8881_) );
AOI21X1 AOI21X1_504 ( .A(_7624__bF_buf2), .B(_8877_), .C(_8881_), .Y(_8882_) );
NAND2X1 NAND2X1_540 ( .A(_6638_), .B(_7569__bF_buf9), .Y(_8883_) );
OAI21X1 OAI21X1_1710 ( .A(cpuregs_29_[17]), .B(_7569__bF_buf8), .C(_8883_), .Y(_8884_) );
NAND2X1 NAND2X1_541 ( .A(decoded_rs1_0_bF_buf3_), .B(_6641_), .Y(_8885_) );
OAI21X1 OAI21X1_1711 ( .A(cpuregs_30_[17]), .B(decoded_rs1_0_bF_buf2_), .C(_8885_), .Y(_8886_) );
MUX2X1 MUX2X1_171 ( .A(_8884_), .B(_8886_), .S(_7556__bF_buf16), .Y(_8887_) );
AND2X2 AND2X2_97 ( .A(cpuregs_25_[17]), .B(decoded_rs1_0_bF_buf1_), .Y(_8888_) );
OAI21X1 OAI21X1_1712 ( .A(_6645_), .B(decoded_rs1_0_bF_buf0_), .C(_7556__bF_buf15), .Y(_8889_) );
AND2X2 AND2X2_98 ( .A(_7569__bF_buf7), .B(cpuregs_26_[17]), .Y(_8890_) );
OAI21X1 OAI21X1_1713 ( .A(_6648_), .B(_7569__bF_buf6), .C(decoded_rs1_1_bF_buf18_), .Y(_8891_) );
OAI22X1 OAI22X1_168 ( .A(_8889_), .B(_8888_), .C(_8891_), .D(_8890_), .Y(_8892_) );
OAI21X1 OAI21X1_1714 ( .A(_8892_), .B(decoded_rs1_2_bF_buf4_), .C(decoded_rs1_3_bF_buf2_), .Y(_8893_) );
AOI21X1 AOI21X1_505 ( .A(decoded_rs1_2_bF_buf3_), .B(_8887_), .C(_8893_), .Y(_8894_) );
AOI21X1 AOI21X1_506 ( .A(decoded_rs1_2_bF_buf2_), .B(_6610_), .C(_7569__bF_buf5), .Y(_8895_) );
OAI21X1 OAI21X1_1715 ( .A(cpuregs_17_[17]), .B(decoded_rs1_2_bF_buf1_), .C(_8895_), .Y(_8896_) );
AOI21X1 AOI21X1_507 ( .A(decoded_rs1_2_bF_buf0_), .B(_6607_), .C(decoded_rs1_0_bF_buf57_), .Y(_8897_) );
OAI21X1 OAI21X1_1716 ( .A(cpuregs_16_[17]), .B(decoded_rs1_2_bF_buf12_), .C(_8897_), .Y(_8898_) );
NAND3X1 NAND3X1_40 ( .A(_7556__bF_buf14), .B(_8896_), .C(_8898_), .Y(_8899_) );
AOI21X1 AOI21X1_508 ( .A(decoded_rs1_2_bF_buf11_), .B(_6617_), .C(_7569__bF_buf4), .Y(_8900_) );
OAI21X1 OAI21X1_1717 ( .A(cpuregs_19_[17]), .B(decoded_rs1_2_bF_buf10_), .C(_8900_), .Y(_8901_) );
AOI21X1 AOI21X1_509 ( .A(decoded_rs1_2_bF_buf9_), .B(_6614_), .C(decoded_rs1_0_bF_buf56_), .Y(_8902_) );
OAI21X1 OAI21X1_1718 ( .A(cpuregs_18_[17]), .B(decoded_rs1_2_bF_buf8_), .C(_8902_), .Y(_8903_) );
NAND3X1 NAND3X1_41 ( .A(decoded_rs1_1_bF_buf17_), .B(_8901_), .C(_8903_), .Y(_8904_) );
AOI21X1 AOI21X1_510 ( .A(_8899_), .B(_8904_), .C(decoded_rs1_3_bF_buf1_), .Y(_8905_) );
OAI21X1 OAI21X1_1719 ( .A(_8894_), .B(_8905_), .C(decoded_rs1_4_bF_buf1_), .Y(_8906_) );
NOR2X1 NOR2X1_735 ( .A(_6653_), .B(_7569__bF_buf3), .Y(_8907_) );
OAI21X1 OAI21X1_1720 ( .A(_6657_), .B(decoded_rs1_0_bF_buf55_), .C(_7556__bF_buf13), .Y(_8908_) );
INVX1 INVX1_735 ( .A(cpuregs_10_[17]), .Y(_8909_) );
AOI21X1 AOI21X1_511 ( .A(cpuregs_11_[17]), .B(decoded_rs1_0_bF_buf54_), .C(_7556__bF_buf12), .Y(_8910_) );
OAI21X1 OAI21X1_1721 ( .A(_8909_), .B(decoded_rs1_0_bF_buf53_), .C(_8910_), .Y(_8911_) );
OAI21X1 OAI21X1_1722 ( .A(_8907_), .B(_8908_), .C(_8911_), .Y(_8912_) );
NOR2X1 NOR2X1_736 ( .A(decoded_rs1_2_bF_buf7_), .B(_8912_), .Y(_8913_) );
NOR2X1 NOR2X1_737 ( .A(_6660_), .B(_7569__bF_buf2), .Y(_8914_) );
OAI21X1 OAI21X1_1723 ( .A(_6664_), .B(decoded_rs1_0_bF_buf52_), .C(_7556__bF_buf11), .Y(_8915_) );
INVX1 INVX1_736 ( .A(cpuregs_14_[17]), .Y(_8916_) );
AOI21X1 AOI21X1_512 ( .A(cpuregs_15_[17]), .B(decoded_rs1_0_bF_buf51_), .C(_7556__bF_buf10), .Y(_8917_) );
OAI21X1 OAI21X1_1724 ( .A(_8916_), .B(decoded_rs1_0_bF_buf50_), .C(_8917_), .Y(_8918_) );
OAI21X1 OAI21X1_1725 ( .A(_8914_), .B(_8915_), .C(_8918_), .Y(_8919_) );
OAI21X1 OAI21X1_1726 ( .A(_8919_), .B(_7560__bF_buf10), .C(decoded_rs1_3_bF_buf0_), .Y(_8920_) );
NAND2X1 NAND2X1_542 ( .A(_6622_), .B(_7569__bF_buf1), .Y(_8921_) );
OAI21X1 OAI21X1_1727 ( .A(cpuregs_1_[17]), .B(_7569__bF_buf0), .C(_8921_), .Y(_8922_) );
NAND2X1 NAND2X1_543 ( .A(_6625_), .B(_7569__bF_buf48), .Y(_8923_) );
OAI21X1 OAI21X1_1728 ( .A(cpuregs_3_[17]), .B(_7569__bF_buf47), .C(_8923_), .Y(_8924_) );
MUX2X1 MUX2X1_172 ( .A(_8924_), .B(_8922_), .S(decoded_rs1_1_bF_buf16_), .Y(_8925_) );
MUX2X1 MUX2X1_173 ( .A(cpuregs_6_[17]), .B(cpuregs_4_[17]), .S(decoded_rs1_1_bF_buf15_), .Y(_8926_) );
NOR2X1 NOR2X1_738 ( .A(decoded_rs1_0_bF_buf49_), .B(_8926_), .Y(_8927_) );
MUX2X1 MUX2X1_174 ( .A(cpuregs_7_[17]), .B(cpuregs_5_[17]), .S(decoded_rs1_1_bF_buf14_), .Y(_8928_) );
OAI21X1 OAI21X1_1729 ( .A(_8928_), .B(_7569__bF_buf46), .C(decoded_rs1_2_bF_buf6_), .Y(_8929_) );
OAI22X1 OAI22X1_169 ( .A(_8927_), .B(_8929_), .C(_8925_), .D(decoded_rs1_2_bF_buf5_), .Y(_8930_) );
NAND2X1 NAND2X1_544 ( .A(_7561__bF_buf6), .B(_8930_), .Y(_8931_) );
OAI21X1 OAI21X1_1730 ( .A(_8913_), .B(_8920_), .C(_8931_), .Y(_8932_) );
AOI21X1 AOI21X1_513 ( .A(_7552__bF_buf5), .B(_8932_), .C(_7586__bF_buf2), .Y(_8933_) );
AOI22X1 AOI22X1_78 ( .A(reg_pc_17_), .B(_7551__bF_buf2), .C(_8933_), .D(_8906_), .Y(_8934_) );
OAI21X1 OAI21X1_1731 ( .A(_4597__bF_buf0), .B(_8855_), .C(_10734__17_), .Y(_8935_) );
OAI21X1 OAI21X1_1732 ( .A(_8934_), .B(_4538__bF_buf2), .C(_8935_), .Y(_8936_) );
NOR2X1 NOR2X1_739 ( .A(_8936_), .B(_8882_), .Y(_8937_) );
AND2X2 AND2X2_99 ( .A(_8937_), .B(_8880_), .Y(_8938_) );
NOR2X1 NOR2X1_740 ( .A(_5217_), .B(_7698__bF_buf3), .Y(_8939_) );
OAI21X1 OAI21X1_1733 ( .A(_5196_), .B(_7700__bF_buf2), .C(_4580__bF_buf4), .Y(_8940_) );
OAI21X1 OAI21X1_1734 ( .A(_5051_), .B(_7700__bF_buf1), .C(_4579__bF_buf1), .Y(_8941_) );
OAI22X1 OAI22X1_170 ( .A(_8694_), .B(_8941_), .C(_8940_), .D(_8939_), .Y(_8942_) );
NOR2X1 NOR2X1_741 ( .A(_8942_), .B(_7697__bF_buf0), .Y(_8943_) );
NOR2X1 NOR2X1_742 ( .A(_4426__bF_buf2), .B(_8943_), .Y(_8944_) );
AOI22X1 AOI22X1_79 ( .A(_4426__bF_buf1), .B(_5057_), .C(_8938_), .D(_8944_), .Y(_81__17_) );
NOR2X1 NOR2X1_743 ( .A(_8869_), .B(_8876_), .Y(_8945_) );
NAND2X1 NAND2X1_545 ( .A(_10734__18_), .B(decoded_imm_18_), .Y(_8946_) );
INVX1 INVX1_737 ( .A(decoded_imm_18_), .Y(_8947_) );
NAND2X1 NAND2X1_546 ( .A(_5045_), .B(_8947_), .Y(_8948_) );
NAND2X1 NAND2X1_547 ( .A(_8946_), .B(_8948_), .Y(_8949_) );
XNOR2X1 XNOR2X1_10 ( .A(_8945_), .B(_8949_), .Y(_8950_) );
NAND2X1 NAND2X1_548 ( .A(_7632__bF_buf3), .B(_8950_), .Y(_8951_) );
AOI21X1 AOI21X1_514 ( .A(_5045_), .B(_7631__bF_buf1), .C(_7629__bF_buf3), .Y(_8952_) );
NAND2X1 NAND2X1_549 ( .A(_8952_), .B(_8951_), .Y(_8953_) );
OAI21X1 OAI21X1_1735 ( .A(_7624__bF_buf1), .B(_10734__18_), .C(cpu_state_5_bF_buf1_), .Y(_8954_) );
AOI21X1 AOI21X1_515 ( .A(_7624__bF_buf0), .B(_8950_), .C(_8954_), .Y(_8955_) );
AND2X2 AND2X2_100 ( .A(cpuregs_17_[18]), .B(decoded_rs1_0_bF_buf48_), .Y(_8956_) );
INVX1 INVX1_738 ( .A(cpuregs_16_[18]), .Y(_8957_) );
OAI21X1 OAI21X1_1736 ( .A(_8957_), .B(decoded_rs1_0_bF_buf47_), .C(_7556__bF_buf9), .Y(_8958_) );
AND2X2 AND2X2_101 ( .A(_7569__bF_buf45), .B(cpuregs_18_[18]), .Y(_8959_) );
INVX1 INVX1_739 ( .A(cpuregs_19_[18]), .Y(_8960_) );
OAI21X1 OAI21X1_1737 ( .A(_8960_), .B(_7569__bF_buf44), .C(decoded_rs1_1_bF_buf13_), .Y(_8961_) );
OAI22X1 OAI22X1_171 ( .A(_8958_), .B(_8956_), .C(_8961_), .D(_8959_), .Y(_8962_) );
NOR2X1 NOR2X1_744 ( .A(decoded_rs1_2_bF_buf4_), .B(_8962_), .Y(_8963_) );
NOR2X1 NOR2X1_745 ( .A(_6675_), .B(_7569__bF_buf43), .Y(_8964_) );
OAI21X1 OAI21X1_1738 ( .A(_6672_), .B(decoded_rs1_0_bF_buf46_), .C(_7556__bF_buf8), .Y(_8965_) );
NOR2X1 NOR2X1_746 ( .A(decoded_rs1_0_bF_buf45_), .B(_6679_), .Y(_8966_) );
OAI21X1 OAI21X1_1739 ( .A(_6682_), .B(_7569__bF_buf42), .C(decoded_rs1_1_bF_buf12_), .Y(_8967_) );
OAI22X1 OAI22X1_172 ( .A(_8965_), .B(_8964_), .C(_8967_), .D(_8966_), .Y(_8968_) );
OAI21X1 OAI21X1_1740 ( .A(_8968_), .B(_7560__bF_buf9), .C(_7561__bF_buf5), .Y(_8969_) );
NOR2X1 NOR2X1_747 ( .A(_8963_), .B(_8969_), .Y(_8970_) );
AOI21X1 AOI21X1_516 ( .A(_6702_), .B(_7556__bF_buf7), .C(decoded_rs1_0_bF_buf44_), .Y(_8971_) );
OAI21X1 OAI21X1_1741 ( .A(cpuregs_30_[18]), .B(_7556__bF_buf6), .C(_8971_), .Y(_8972_) );
NOR2X1 NOR2X1_748 ( .A(cpuregs_31_[18]), .B(_7556__bF_buf5), .Y(_8973_) );
OAI21X1 OAI21X1_1742 ( .A(cpuregs_29_[18]), .B(decoded_rs1_1_bF_buf11_), .C(decoded_rs1_0_bF_buf43_), .Y(_8974_) );
OAI21X1 OAI21X1_1743 ( .A(_8973_), .B(_8974_), .C(_8972_), .Y(_8975_) );
INVX1 INVX1_740 ( .A(cpuregs_26_[18]), .Y(_8976_) );
OAI21X1 OAI21X1_1744 ( .A(cpuregs_24_[18]), .B(decoded_rs1_1_bF_buf10_), .C(_7569__bF_buf41), .Y(_8977_) );
AOI21X1 AOI21X1_517 ( .A(_8976_), .B(decoded_rs1_1_bF_buf9_), .C(_8977_), .Y(_8978_) );
OAI21X1 OAI21X1_1745 ( .A(cpuregs_25_[18]), .B(decoded_rs1_1_bF_buf8_), .C(decoded_rs1_0_bF_buf42_), .Y(_8979_) );
AOI21X1 AOI21X1_518 ( .A(_6713_), .B(decoded_rs1_1_bF_buf7_), .C(_8979_), .Y(_8980_) );
OAI21X1 OAI21X1_1746 ( .A(_8978_), .B(_8980_), .C(_7560__bF_buf8), .Y(_8981_) );
NAND2X1 NAND2X1_550 ( .A(decoded_rs1_3_bF_buf6_), .B(_8981_), .Y(_8982_) );
AOI21X1 AOI21X1_519 ( .A(decoded_rs1_2_bF_buf3_), .B(_8975_), .C(_8982_), .Y(_8983_) );
OAI21X1 OAI21X1_1747 ( .A(_8983_), .B(_8970_), .C(decoded_rs1_4_bF_buf0_), .Y(_8984_) );
INVX1 INVX1_741 ( .A(cpuregs_14_[18]), .Y(_8985_) );
OAI21X1 OAI21X1_1748 ( .A(cpuregs_12_[18]), .B(decoded_rs1_1_bF_buf6_), .C(_7569__bF_buf40), .Y(_8986_) );
AOI21X1 AOI21X1_520 ( .A(_8985_), .B(decoded_rs1_1_bF_buf5_), .C(_8986_), .Y(_8987_) );
INVX1 INVX1_742 ( .A(cpuregs_15_[18]), .Y(_8988_) );
OAI21X1 OAI21X1_1749 ( .A(cpuregs_13_[18]), .B(decoded_rs1_1_bF_buf4_), .C(decoded_rs1_0_bF_buf41_), .Y(_8989_) );
AOI21X1 AOI21X1_521 ( .A(_8988_), .B(decoded_rs1_1_bF_buf3_), .C(_8989_), .Y(_8990_) );
OAI21X1 OAI21X1_1750 ( .A(_8987_), .B(_8990_), .C(decoded_rs1_2_bF_buf2_), .Y(_8991_) );
INVX1 INVX1_743 ( .A(cpuregs_10_[18]), .Y(_8992_) );
OAI21X1 OAI21X1_1751 ( .A(cpuregs_8_[18]), .B(decoded_rs1_1_bF_buf2_), .C(_7569__bF_buf39), .Y(_8993_) );
AOI21X1 AOI21X1_522 ( .A(_8992_), .B(decoded_rs1_1_bF_buf1_), .C(_8993_), .Y(_8994_) );
INVX1 INVX1_744 ( .A(cpuregs_11_[18]), .Y(_8995_) );
OAI21X1 OAI21X1_1752 ( .A(cpuregs_9_[18]), .B(decoded_rs1_1_bF_buf0_), .C(decoded_rs1_0_bF_buf40_), .Y(_8996_) );
AOI21X1 AOI21X1_523 ( .A(_8995_), .B(decoded_rs1_1_bF_buf44_), .C(_8996_), .Y(_8997_) );
OAI21X1 OAI21X1_1753 ( .A(_8994_), .B(_8997_), .C(_7560__bF_buf7), .Y(_8998_) );
NAND2X1 NAND2X1_551 ( .A(_8998_), .B(_8991_), .Y(_8999_) );
AND2X2 AND2X2_102 ( .A(cpuregs_1_[18]), .B(decoded_rs1_0_bF_buf39_), .Y(_9000_) );
INVX1 INVX1_745 ( .A(cpuregs_0_[18]), .Y(_9001_) );
OAI21X1 OAI21X1_1754 ( .A(_9001_), .B(decoded_rs1_0_bF_buf38_), .C(_7556__bF_buf4), .Y(_9002_) );
NOR2X1 NOR2X1_749 ( .A(decoded_rs1_0_bF_buf37_), .B(_6693_), .Y(_9003_) );
INVX1 INVX1_746 ( .A(cpuregs_3_[18]), .Y(_9004_) );
OAI21X1 OAI21X1_1755 ( .A(_9004_), .B(_7569__bF_buf38), .C(decoded_rs1_1_bF_buf43_), .Y(_9005_) );
OAI22X1 OAI22X1_173 ( .A(_9002_), .B(_9000_), .C(_9005_), .D(_9003_), .Y(_9006_) );
NOR2X1 NOR2X1_750 ( .A(decoded_rs1_2_bF_buf1_), .B(_9006_), .Y(_9007_) );
AND2X2 AND2X2_103 ( .A(cpuregs_5_[18]), .B(decoded_rs1_0_bF_buf36_), .Y(_9008_) );
INVX1 INVX1_747 ( .A(cpuregs_4_[18]), .Y(_9009_) );
OAI21X1 OAI21X1_1756 ( .A(_9009_), .B(decoded_rs1_0_bF_buf35_), .C(_7556__bF_buf3), .Y(_9010_) );
NOR2X1 NOR2X1_751 ( .A(decoded_rs1_0_bF_buf34_), .B(_6687_), .Y(_9011_) );
INVX1 INVX1_748 ( .A(cpuregs_7_[18]), .Y(_9012_) );
OAI21X1 OAI21X1_1757 ( .A(_9012_), .B(_7569__bF_buf37), .C(decoded_rs1_1_bF_buf42_), .Y(_9013_) );
OAI22X1 OAI22X1_174 ( .A(_9010_), .B(_9008_), .C(_9013_), .D(_9011_), .Y(_9014_) );
OAI21X1 OAI21X1_1758 ( .A(_9014_), .B(_7560__bF_buf6), .C(_7561__bF_buf4), .Y(_9015_) );
OAI22X1 OAI22X1_175 ( .A(_9007_), .B(_9015_), .C(_8999_), .D(_7561__bF_buf3), .Y(_9016_) );
AOI21X1 AOI21X1_524 ( .A(_7552__bF_buf4), .B(_9016_), .C(_7586__bF_buf1), .Y(_9017_) );
AOI22X1 AOI22X1_80 ( .A(reg_pc_18_), .B(_7551__bF_buf1), .C(_9017_), .D(_8984_), .Y(_9018_) );
OAI21X1 OAI21X1_1759 ( .A(instr_slli), .B(instr_sll), .C(_10734__17_), .Y(_9019_) );
OAI21X1 OAI21X1_1760 ( .A(_7698__bF_buf2), .B(_5040_), .C(_9019_), .Y(_9020_) );
INVX1 INVX1_749 ( .A(_10734__22_), .Y(_9021_) );
OAI21X1 OAI21X1_1761 ( .A(_7698__bF_buf1), .B(_9021_), .C(_8764_), .Y(_9022_) );
MUX2X1 MUX2X1_175 ( .A(_9020_), .B(_9022_), .S(_4579__bF_buf0), .Y(_9023_) );
OR2X2 OR2X2_9 ( .A(_7697__bF_buf3), .B(_9023_), .Y(_9024_) );
OAI21X1 OAI21X1_1762 ( .A(_7627_), .B(_5045_), .C(resetn_bF_buf5), .Y(_9025_) );
AOI21X1 AOI21X1_525 ( .A(_10734__18_), .B(_4597__bF_buf3), .C(_9025_), .Y(_9026_) );
AND2X2 AND2X2_104 ( .A(_9024_), .B(_9026_), .Y(_9027_) );
OAI21X1 OAI21X1_1763 ( .A(_9018_), .B(_4538__bF_buf1), .C(_9027_), .Y(_9028_) );
NOR2X1 NOR2X1_752 ( .A(_9028_), .B(_8955_), .Y(_9029_) );
AOI22X1 AOI22X1_81 ( .A(_4426__bF_buf0), .B(_5045_), .C(_9029_), .D(_8953_), .Y(_81__18_) );
OAI21X1 OAI21X1_1764 ( .A(_8945_), .B(_8949_), .C(_8946_), .Y(_9030_) );
NAND2X1 NAND2X1_552 ( .A(_10734__19_), .B(decoded_imm_19_), .Y(_9031_) );
INVX1 INVX1_750 ( .A(_9031_), .Y(_9032_) );
NOR2X1 NOR2X1_753 ( .A(_10734__19_), .B(decoded_imm_19_), .Y(_9033_) );
OR2X2 OR2X2_10 ( .A(_9032_), .B(_9033_), .Y(_9034_) );
XNOR2X1 XNOR2X1_11 ( .A(_9030_), .B(_9034_), .Y(_9035_) );
AOI21X1 AOI21X1_526 ( .A(_5040_), .B(_7631__bF_buf0), .C(_7629__bF_buf2), .Y(_9036_) );
OAI21X1 OAI21X1_1765 ( .A(_9035_), .B(_7631__bF_buf5), .C(_9036_), .Y(_9037_) );
AOI21X1 AOI21X1_527 ( .A(_5040_), .B(_7623__bF_buf2), .C(_4587__bF_buf1), .Y(_9038_) );
OAI21X1 OAI21X1_1766 ( .A(_9035_), .B(_7623__bF_buf1), .C(_9038_), .Y(_9039_) );
MUX2X1 MUX2X1_176 ( .A(cpuregs_9_[19]), .B(cpuregs_8_[19]), .S(decoded_rs1_0_bF_buf33_), .Y(_9040_) );
MUX2X1 MUX2X1_177 ( .A(cpuregs_11_[19]), .B(cpuregs_10_[19]), .S(decoded_rs1_0_bF_buf32_), .Y(_9041_) );
MUX2X1 MUX2X1_178 ( .A(_9041_), .B(_9040_), .S(decoded_rs1_1_bF_buf41_), .Y(_9042_) );
NOR2X1 NOR2X1_754 ( .A(_6755_), .B(_7569__bF_buf36), .Y(_9043_) );
INVX1 INVX1_751 ( .A(cpuregs_12_[19]), .Y(_9044_) );
OAI21X1 OAI21X1_1767 ( .A(_9044_), .B(decoded_rs1_0_bF_buf31_), .C(_7556__bF_buf2), .Y(_9045_) );
INVX1 INVX1_752 ( .A(cpuregs_14_[19]), .Y(_9046_) );
AOI21X1 AOI21X1_528 ( .A(cpuregs_15_[19]), .B(decoded_rs1_0_bF_buf30_), .C(_7556__bF_buf1), .Y(_9047_) );
OAI21X1 OAI21X1_1768 ( .A(_9046_), .B(decoded_rs1_0_bF_buf29_), .C(_9047_), .Y(_9048_) );
OAI21X1 OAI21X1_1769 ( .A(_9043_), .B(_9045_), .C(_9048_), .Y(_9049_) );
OAI21X1 OAI21X1_1770 ( .A(_9049_), .B(_7560__bF_buf5), .C(decoded_rs1_3_bF_buf5_), .Y(_9050_) );
AOI21X1 AOI21X1_529 ( .A(_7560__bF_buf4), .B(_9042_), .C(_9050_), .Y(_9051_) );
MUX2X1 MUX2X1_179 ( .A(cpuregs_2_[19]), .B(cpuregs_0_[19]), .S(decoded_rs1_1_bF_buf40_), .Y(_9052_) );
NOR2X1 NOR2X1_755 ( .A(decoded_rs1_0_bF_buf28_), .B(_9052_), .Y(_9053_) );
MUX2X1 MUX2X1_180 ( .A(cpuregs_3_[19]), .B(cpuregs_1_[19]), .S(decoded_rs1_1_bF_buf39_), .Y(_9054_) );
OAI21X1 OAI21X1_1771 ( .A(_9054_), .B(_7569__bF_buf35), .C(_7560__bF_buf3), .Y(_9055_) );
MUX2X1 MUX2X1_181 ( .A(cpuregs_6_[19]), .B(cpuregs_4_[19]), .S(decoded_rs1_1_bF_buf38_), .Y(_9056_) );
NOR2X1 NOR2X1_756 ( .A(decoded_rs1_0_bF_buf27_), .B(_9056_), .Y(_9057_) );
MUX2X1 MUX2X1_182 ( .A(cpuregs_7_[19]), .B(cpuregs_5_[19]), .S(decoded_rs1_1_bF_buf37_), .Y(_9058_) );
OAI21X1 OAI21X1_1772 ( .A(_9058_), .B(_7569__bF_buf34), .C(decoded_rs1_2_bF_buf0_), .Y(_9059_) );
OAI22X1 OAI22X1_176 ( .A(_9055_), .B(_9053_), .C(_9057_), .D(_9059_), .Y(_9060_) );
AND2X2 AND2X2_105 ( .A(_9060_), .B(_7561__bF_buf2), .Y(_9061_) );
OAI21X1 OAI21X1_1773 ( .A(_9051_), .B(_9061_), .C(_7552__bF_buf3), .Y(_9062_) );
NOR2X1 NOR2X1_757 ( .A(_6738_), .B(_7569__bF_buf33), .Y(_9063_) );
OAI21X1 OAI21X1_1774 ( .A(_6735_), .B(decoded_rs1_0_bF_buf26_), .C(_7556__bF_buf0), .Y(_9064_) );
NOR2X1 NOR2X1_758 ( .A(decoded_rs1_0_bF_buf25_), .B(_6742_), .Y(_9065_) );
OAI21X1 OAI21X1_1775 ( .A(_6745_), .B(_7569__bF_buf32), .C(decoded_rs1_1_bF_buf36_), .Y(_9066_) );
OAI22X1 OAI22X1_177 ( .A(_9064_), .B(_9063_), .C(_9066_), .D(_9065_), .Y(_9067_) );
MUX2X1 MUX2X1_183 ( .A(cpuregs_25_[19]), .B(cpuregs_24_[19]), .S(decoded_rs1_0_bF_buf24_), .Y(_9068_) );
MUX2X1 MUX2X1_184 ( .A(cpuregs_27_[19]), .B(cpuregs_26_[19]), .S(decoded_rs1_0_bF_buf23_), .Y(_9069_) );
MUX2X1 MUX2X1_185 ( .A(_9068_), .B(_9069_), .S(_7556__bF_buf42), .Y(_9070_) );
AOI21X1 AOI21X1_530 ( .A(_7560__bF_buf2), .B(_9070_), .C(_7561__bF_buf1), .Y(_9071_) );
OAI21X1 OAI21X1_1776 ( .A(_7560__bF_buf1), .B(_9067_), .C(_9071_), .Y(_9072_) );
AOI21X1 AOI21X1_531 ( .A(cpuregs_16_[19]), .B(_7569__bF_buf31), .C(decoded_rs1_1_bF_buf35_), .Y(_9073_) );
OAI21X1 OAI21X1_1777 ( .A(_6764_), .B(_7569__bF_buf30), .C(_9073_), .Y(_9074_) );
AND2X2 AND2X2_106 ( .A(_7569__bF_buf29), .B(cpuregs_18_[19]), .Y(_9075_) );
INVX1 INVX1_753 ( .A(cpuregs_19_[19]), .Y(_9076_) );
OAI21X1 OAI21X1_1778 ( .A(_9076_), .B(_7569__bF_buf28), .C(decoded_rs1_1_bF_buf34_), .Y(_9077_) );
OAI21X1 OAI21X1_1779 ( .A(_9075_), .B(_9077_), .C(_9074_), .Y(_9078_) );
NOR2X1 NOR2X1_759 ( .A(decoded_rs1_2_bF_buf12_), .B(_9078_), .Y(_9079_) );
AND2X2 AND2X2_107 ( .A(cpuregs_21_[19]), .B(decoded_rs1_0_bF_buf22_), .Y(_9080_) );
OAI21X1 OAI21X1_1780 ( .A(_6770_), .B(decoded_rs1_0_bF_buf21_), .C(_7556__bF_buf41), .Y(_9081_) );
AOI21X1 AOI21X1_532 ( .A(cpuregs_23_[19]), .B(decoded_rs1_0_bF_buf20_), .C(_7556__bF_buf40), .Y(_9082_) );
OAI21X1 OAI21X1_1781 ( .A(_6773_), .B(decoded_rs1_0_bF_buf19_), .C(_9082_), .Y(_9083_) );
OAI21X1 OAI21X1_1782 ( .A(_9080_), .B(_9081_), .C(_9083_), .Y(_9084_) );
OAI21X1 OAI21X1_1783 ( .A(_9084_), .B(_7560__bF_buf0), .C(_7561__bF_buf0), .Y(_9085_) );
OAI21X1 OAI21X1_1784 ( .A(_9079_), .B(_9085_), .C(_9072_), .Y(_9086_) );
AOI21X1 AOI21X1_533 ( .A(decoded_rs1_4_bF_buf4_), .B(_9086_), .C(_7586__bF_buf0), .Y(_9087_) );
AOI22X1 AOI22X1_82 ( .A(reg_pc_19_), .B(_7551__bF_buf0), .C(_9087_), .D(_9062_), .Y(_9088_) );
NOR2X1 NOR2X1_760 ( .A(_4538__bF_buf0), .B(_9088_), .Y(_9089_) );
INVX1 INVX1_754 ( .A(_8860_), .Y(_9090_) );
INVX1 INVX1_755 ( .A(_10734__23_), .Y(_9091_) );
OAI21X1 OAI21X1_1785 ( .A(_7698__bF_buf0), .B(_9091_), .C(_4580__bF_buf3), .Y(_9092_) );
OAI21X1 OAI21X1_1786 ( .A(_5045_), .B(_7700__bF_buf0), .C(_4579__bF_buf4), .Y(_9093_) );
OAI22X1 OAI22X1_178 ( .A(_8864_), .B(_9093_), .C(_9092_), .D(_9090_), .Y(_9094_) );
OAI21X1 OAI21X1_1787 ( .A(_7627_), .B(_5040_), .C(resetn_bF_buf4), .Y(_9095_) );
AOI21X1 AOI21X1_534 ( .A(_10734__19_), .B(_4597__bF_buf2), .C(_9095_), .Y(_9096_) );
OAI21X1 OAI21X1_1788 ( .A(_7697__bF_buf2), .B(_9094_), .C(_9096_), .Y(_9097_) );
NOR2X1 NOR2X1_761 ( .A(_9097_), .B(_9089_), .Y(_9098_) );
AND2X2 AND2X2_108 ( .A(_9039_), .B(_9098_), .Y(_9099_) );
AOI22X1 AOI22X1_83 ( .A(_4426__bF_buf11), .B(_5040_), .C(_9099_), .D(_9037_), .Y(_81__19_) );
OAI21X1 OAI21X1_1789 ( .A(_5057_), .B(_8868_), .C(_8874_), .Y(_9100_) );
NOR2X1 NOR2X1_762 ( .A(_8949_), .B(_9034_), .Y(_9101_) );
OAI21X1 OAI21X1_1790 ( .A(_9033_), .B(_8946_), .C(_9031_), .Y(_9102_) );
AOI21X1 AOI21X1_535 ( .A(_9101_), .B(_9100_), .C(_9102_), .Y(_9103_) );
INVX1 INVX1_756 ( .A(_9101_), .Y(_9104_) );
OR2X2 OR2X2_11 ( .A(_9104_), .B(_8875_), .Y(_9105_) );
OAI21X1 OAI21X1_1791 ( .A(_8781_), .B(_9105_), .C(_9103_), .Y(_9106_) );
INVX1 INVX1_757 ( .A(decoded_imm_20_), .Y(_9107_) );
NAND2X1 NAND2X1_553 ( .A(_5218_), .B(_9107_), .Y(_9108_) );
NAND2X1 NAND2X1_554 ( .A(_10734__20_), .B(decoded_imm_20_), .Y(_9109_) );
NAND2X1 NAND2X1_555 ( .A(_9109_), .B(_9108_), .Y(_9110_) );
INVX1 INVX1_758 ( .A(_9110_), .Y(_9111_) );
XNOR2X1 XNOR2X1_12 ( .A(_9106_), .B(_9111_), .Y(_9112_) );
OAI21X1 OAI21X1_1792 ( .A(_7632__bF_buf2), .B(_10734__20_), .C(_7630_), .Y(_9113_) );
AOI21X1 AOI21X1_536 ( .A(_7632__bF_buf1), .B(_9112_), .C(_9113_), .Y(_9114_) );
OAI21X1 OAI21X1_1793 ( .A(_7624__bF_buf4), .B(_10734__20_), .C(cpu_state_5_bF_buf0_), .Y(_9115_) );
AOI21X1 AOI21X1_537 ( .A(_7624__bF_buf3), .B(_9112_), .C(_9115_), .Y(_9116_) );
NOR2X1 NOR2X1_763 ( .A(_6807_), .B(_7569__bF_buf27), .Y(_9117_) );
INVX1 INVX1_759 ( .A(cpuregs_16_[20]), .Y(_9118_) );
OAI21X1 OAI21X1_1794 ( .A(_9118_), .B(decoded_rs1_0_bF_buf18_), .C(_7556__bF_buf39), .Y(_9119_) );
NOR2X1 NOR2X1_764 ( .A(decoded_rs1_0_bF_buf17_), .B(_6810_), .Y(_9120_) );
INVX1 INVX1_760 ( .A(cpuregs_19_[20]), .Y(_9121_) );
OAI21X1 OAI21X1_1795 ( .A(_9121_), .B(_7569__bF_buf26), .C(decoded_rs1_1_bF_buf33_), .Y(_9122_) );
OAI22X1 OAI22X1_179 ( .A(_9119_), .B(_9117_), .C(_9122_), .D(_9120_), .Y(_9123_) );
NOR2X1 NOR2X1_765 ( .A(decoded_rs1_2_bF_buf11_), .B(_9123_), .Y(_9124_) );
NOR2X1 NOR2X1_766 ( .A(_6814_), .B(_7569__bF_buf25), .Y(_9125_) );
INVX1 INVX1_761 ( .A(cpuregs_20_[20]), .Y(_9126_) );
OAI21X1 OAI21X1_1796 ( .A(_9126_), .B(decoded_rs1_0_bF_buf16_), .C(_7556__bF_buf38), .Y(_9127_) );
AND2X2 AND2X2_109 ( .A(_7569__bF_buf24), .B(cpuregs_22_[20]), .Y(_9128_) );
INVX1 INVX1_762 ( .A(cpuregs_23_[20]), .Y(_9129_) );
OAI21X1 OAI21X1_1797 ( .A(_9129_), .B(_7569__bF_buf23), .C(decoded_rs1_1_bF_buf32_), .Y(_9130_) );
OAI22X1 OAI22X1_180 ( .A(_9127_), .B(_9125_), .C(_9130_), .D(_9128_), .Y(_9131_) );
OAI21X1 OAI21X1_1798 ( .A(_9131_), .B(_7560__bF_buf12), .C(_7561__bF_buf6), .Y(_9132_) );
NOR2X1 NOR2X1_767 ( .A(_9124_), .B(_9132_), .Y(_9133_) );
AOI21X1 AOI21X1_538 ( .A(_6795_), .B(_7556__bF_buf37), .C(decoded_rs1_0_bF_buf15_), .Y(_9134_) );
OAI21X1 OAI21X1_1799 ( .A(cpuregs_26_[20]), .B(_7556__bF_buf36), .C(_9134_), .Y(_9135_) );
NOR2X1 NOR2X1_768 ( .A(cpuregs_27_[20]), .B(_7556__bF_buf35), .Y(_9136_) );
OAI21X1 OAI21X1_1800 ( .A(cpuregs_25_[20]), .B(decoded_rs1_1_bF_buf31_), .C(decoded_rs1_0_bF_buf14_), .Y(_9137_) );
OAI21X1 OAI21X1_1801 ( .A(_9136_), .B(_9137_), .C(_9135_), .Y(_9138_) );
NOR2X1 NOR2X1_769 ( .A(cpuregs_30_[20]), .B(_7556__bF_buf34), .Y(_9139_) );
OAI21X1 OAI21X1_1802 ( .A(cpuregs_28_[20]), .B(decoded_rs1_1_bF_buf30_), .C(_7569__bF_buf22), .Y(_9140_) );
NOR2X1 NOR2X1_770 ( .A(cpuregs_31_[20]), .B(_7556__bF_buf33), .Y(_9141_) );
OAI21X1 OAI21X1_1803 ( .A(cpuregs_29_[20]), .B(decoded_rs1_1_bF_buf29_), .C(decoded_rs1_0_bF_buf13_), .Y(_9142_) );
OAI22X1 OAI22X1_181 ( .A(_9139_), .B(_9140_), .C(_9141_), .D(_9142_), .Y(_9143_) );
NAND2X1 NAND2X1_556 ( .A(decoded_rs1_2_bF_buf10_), .B(_9143_), .Y(_9144_) );
NAND2X1 NAND2X1_557 ( .A(decoded_rs1_3_bF_buf4_), .B(_9144_), .Y(_9145_) );
AOI21X1 AOI21X1_539 ( .A(_7560__bF_buf11), .B(_9138_), .C(_9145_), .Y(_9146_) );
OAI21X1 OAI21X1_1804 ( .A(_9146_), .B(_9133_), .C(decoded_rs1_4_bF_buf3_), .Y(_9147_) );
AOI21X1 AOI21X1_540 ( .A(_6830_), .B(_7556__bF_buf32), .C(decoded_rs1_0_bF_buf12_), .Y(_9148_) );
OAI21X1 OAI21X1_1805 ( .A(cpuregs_14_[20]), .B(_7556__bF_buf31), .C(_9148_), .Y(_9149_) );
INVX1 INVX1_763 ( .A(cpuregs_13_[20]), .Y(_9150_) );
AOI21X1 AOI21X1_541 ( .A(_9150_), .B(_7556__bF_buf30), .C(_7569__bF_buf21), .Y(_9151_) );
OAI21X1 OAI21X1_1806 ( .A(cpuregs_15_[20]), .B(_7556__bF_buf29), .C(_9151_), .Y(_9152_) );
AOI21X1 AOI21X1_542 ( .A(_9149_), .B(_9152_), .C(_7560__bF_buf10), .Y(_9153_) );
AND2X2 AND2X2_110 ( .A(cpuregs_1_[20]), .B(decoded_rs1_0_bF_buf11_), .Y(_9154_) );
INVX1 INVX1_764 ( .A(cpuregs_0_[20]), .Y(_9155_) );
OAI21X1 OAI21X1_1807 ( .A(_9155_), .B(decoded_rs1_0_bF_buf10_), .C(_7556__bF_buf28), .Y(_9156_) );
AND2X2 AND2X2_111 ( .A(_7569__bF_buf20), .B(cpuregs_2_[20]), .Y(_9157_) );
INVX1 INVX1_765 ( .A(cpuregs_3_[20]), .Y(_9158_) );
OAI21X1 OAI21X1_1808 ( .A(_9158_), .B(_7569__bF_buf19), .C(decoded_rs1_1_bF_buf28_), .Y(_9159_) );
OAI22X1 OAI22X1_182 ( .A(_9156_), .B(_9154_), .C(_9159_), .D(_9157_), .Y(_9160_) );
NOR2X1 NOR2X1_771 ( .A(decoded_rs1_2_bF_buf9_), .B(_9160_), .Y(_9161_) );
AND2X2 AND2X2_112 ( .A(cpuregs_5_[20]), .B(decoded_rs1_0_bF_buf9_), .Y(_9162_) );
OAI21X1 OAI21X1_1809 ( .A(_6844_), .B(decoded_rs1_0_bF_buf8_), .C(_7556__bF_buf27), .Y(_9163_) );
NOR2X1 NOR2X1_772 ( .A(decoded_rs1_0_bF_buf7_), .B(_6847_), .Y(_9164_) );
INVX1 INVX1_766 ( .A(cpuregs_7_[20]), .Y(_9165_) );
OAI21X1 OAI21X1_1810 ( .A(_9165_), .B(_7569__bF_buf18), .C(decoded_rs1_1_bF_buf27_), .Y(_9166_) );
OAI22X1 OAI22X1_183 ( .A(_9163_), .B(_9162_), .C(_9166_), .D(_9164_), .Y(_9167_) );
OAI21X1 OAI21X1_1811 ( .A(_9167_), .B(_7560__bF_buf9), .C(_7561__bF_buf5), .Y(_9168_) );
AND2X2 AND2X2_113 ( .A(cpuregs_9_[20]), .B(decoded_rs1_0_bF_buf6_), .Y(_9169_) );
OAI21X1 OAI21X1_1812 ( .A(_6823_), .B(decoded_rs1_0_bF_buf5_), .C(_7556__bF_buf26), .Y(_9170_) );
AND2X2 AND2X2_114 ( .A(_7569__bF_buf17), .B(cpuregs_10_[20]), .Y(_9171_) );
OAI21X1 OAI21X1_1813 ( .A(_6826_), .B(_7569__bF_buf16), .C(decoded_rs1_1_bF_buf26_), .Y(_9172_) );
OAI22X1 OAI22X1_184 ( .A(_9170_), .B(_9169_), .C(_9172_), .D(_9171_), .Y(_9173_) );
OAI21X1 OAI21X1_1814 ( .A(_9173_), .B(decoded_rs1_2_bF_buf8_), .C(decoded_rs1_3_bF_buf3_), .Y(_9174_) );
OAI22X1 OAI22X1_185 ( .A(_9168_), .B(_9161_), .C(_9153_), .D(_9174_), .Y(_9175_) );
AOI21X1 AOI21X1_543 ( .A(_7552__bF_buf2), .B(_9175_), .C(_7586__bF_buf3), .Y(_9176_) );
AOI22X1 AOI22X1_84 ( .A(reg_pc_20_), .B(_7551__bF_buf3), .C(_9147_), .D(_9176_), .Y(_9177_) );
OAI21X1 OAI21X1_1815 ( .A(_4597__bF_buf1), .B(_8855_), .C(_10734__20_), .Y(_9178_) );
OAI21X1 OAI21X1_1816 ( .A(_9177_), .B(_4538__bF_buf4), .C(_9178_), .Y(_9179_) );
OR2X2 OR2X2_12 ( .A(_9116_), .B(_9179_), .Y(_9180_) );
NOR2X1 NOR2X1_773 ( .A(_9114_), .B(_9180_), .Y(_9181_) );
OAI21X1 OAI21X1_1817 ( .A(instr_slli), .B(instr_sll), .C(_10734__19_), .Y(_9182_) );
INVX1 INVX1_767 ( .A(_9182_), .Y(_9183_) );
OAI21X1 OAI21X1_1818 ( .A(_8939_), .B(_9183_), .C(_4579__bF_buf3), .Y(_9184_) );
AOI22X1 AOI22X1_85 ( .A(_10734__16_), .B(_8139_), .C(_7616_), .D(_10734__24_), .Y(_9185_) );
OAI21X1 OAI21X1_1819 ( .A(_9185_), .B(_4579__bF_buf2), .C(_9184_), .Y(_9186_) );
AOI21X1 AOI21X1_544 ( .A(_9186_), .B(_4584_), .C(_4426__bF_buf10), .Y(_9187_) );
AOI22X1 AOI22X1_86 ( .A(_4426__bF_buf9), .B(_5218_), .C(_9181_), .D(_9187_), .Y(_81__20_) );
NAND2X1 NAND2X1_558 ( .A(_10734__21_), .B(decoded_imm_21_), .Y(_9188_) );
NOR2X1 NOR2X1_774 ( .A(_10734__21_), .B(decoded_imm_21_), .Y(_9189_) );
INVX1 INVX1_768 ( .A(_9189_), .Y(_9190_) );
NAND2X1 NAND2X1_559 ( .A(_9188_), .B(_9190_), .Y(_9191_) );
NAND2X1 NAND2X1_560 ( .A(_9111_), .B(_9106_), .Y(_9192_) );
OAI21X1 OAI21X1_1820 ( .A(_5218_), .B(_9107_), .C(_9192_), .Y(_9193_) );
XOR2X1 XOR2X1_8 ( .A(_9193_), .B(_9191_), .Y(_9194_) );
NAND2X1 NAND2X1_561 ( .A(_7632__bF_buf0), .B(_9194_), .Y(_9195_) );
AOI21X1 AOI21X1_545 ( .A(_5217_), .B(_7631__bF_buf4), .C(_7629__bF_buf1), .Y(_9196_) );
NAND2X1 NAND2X1_562 ( .A(_9196_), .B(_9195_), .Y(_9197_) );
OAI21X1 OAI21X1_1821 ( .A(_7624__bF_buf2), .B(_10734__21_), .C(cpu_state_5_bF_buf3_), .Y(_9198_) );
AOI21X1 AOI21X1_546 ( .A(_7624__bF_buf1), .B(_9194_), .C(_9198_), .Y(_9199_) );
OAI21X1 OAI21X1_1822 ( .A(_6897_), .B(decoded_rs1_0_bF_buf4_), .C(_7556__bF_buf25), .Y(_9200_) );
AOI21X1 AOI21X1_547 ( .A(cpuregs_17_[21]), .B(decoded_rs1_0_bF_buf3_), .C(_9200_), .Y(_9201_) );
OAI21X1 OAI21X1_1823 ( .A(_6900_), .B(_7569__bF_buf15), .C(decoded_rs1_1_bF_buf25_), .Y(_9202_) );
AOI21X1 AOI21X1_548 ( .A(cpuregs_18_[21]), .B(_7569__bF_buf14), .C(_9202_), .Y(_9203_) );
OAI21X1 OAI21X1_1824 ( .A(_9203_), .B(_9201_), .C(_7560__bF_buf8), .Y(_9204_) );
NOR2X1 NOR2X1_775 ( .A(cpuregs_20_[21]), .B(decoded_rs1_0_bF_buf2_), .Y(_9205_) );
AOI21X1 AOI21X1_549 ( .A(_6905_), .B(decoded_rs1_0_bF_buf1_), .C(_9205_), .Y(_9206_) );
AOI21X1 AOI21X1_550 ( .A(cpuregs_23_[21]), .B(decoded_rs1_0_bF_buf0_), .C(_7556__bF_buf24), .Y(_9207_) );
OAI21X1 OAI21X1_1825 ( .A(_6908_), .B(decoded_rs1_0_bF_buf57_), .C(_9207_), .Y(_9208_) );
OAI21X1 OAI21X1_1826 ( .A(decoded_rs1_1_bF_buf24_), .B(_9206_), .C(_9208_), .Y(_9209_) );
NAND2X1 NAND2X1_563 ( .A(decoded_rs1_2_bF_buf7_), .B(_9209_), .Y(_9210_) );
AOI21X1 AOI21X1_551 ( .A(_9204_), .B(_9210_), .C(decoded_rs1_3_bF_buf2_), .Y(_9211_) );
OAI21X1 OAI21X1_1827 ( .A(_6889_), .B(decoded_rs1_0_bF_buf56_), .C(_7556__bF_buf23), .Y(_9212_) );
AOI21X1 AOI21X1_552 ( .A(cpuregs_29_[21]), .B(decoded_rs1_0_bF_buf55_), .C(_9212_), .Y(_9213_) );
INVX1 INVX1_769 ( .A(cpuregs_31_[21]), .Y(_9214_) );
OAI21X1 OAI21X1_1828 ( .A(_9214_), .B(_7569__bF_buf13), .C(decoded_rs1_1_bF_buf23_), .Y(_9215_) );
AOI21X1 AOI21X1_553 ( .A(cpuregs_30_[21]), .B(_7569__bF_buf12), .C(_9215_), .Y(_9216_) );
OAI21X1 OAI21X1_1829 ( .A(_9216_), .B(_9213_), .C(decoded_rs1_2_bF_buf6_), .Y(_9217_) );
OAI21X1 OAI21X1_1830 ( .A(_6886_), .B(decoded_rs1_0_bF_buf54_), .C(_7556__bF_buf22), .Y(_9218_) );
AOI21X1 AOI21X1_554 ( .A(cpuregs_25_[21]), .B(decoded_rs1_0_bF_buf53_), .C(_9218_), .Y(_9219_) );
INVX1 INVX1_770 ( .A(cpuregs_27_[21]), .Y(_9220_) );
OAI21X1 OAI21X1_1831 ( .A(_9220_), .B(_7569__bF_buf11), .C(decoded_rs1_1_bF_buf22_), .Y(_9221_) );
AOI21X1 AOI21X1_555 ( .A(cpuregs_26_[21]), .B(_7569__bF_buf10), .C(_9221_), .Y(_9222_) );
OAI21X1 OAI21X1_1832 ( .A(_9222_), .B(_9219_), .C(_7560__bF_buf7), .Y(_9223_) );
AOI21X1 AOI21X1_556 ( .A(_9217_), .B(_9223_), .C(_7561__bF_buf4), .Y(_9224_) );
OAI21X1 OAI21X1_1833 ( .A(_9211_), .B(_9224_), .C(decoded_rs1_4_bF_buf2_), .Y(_9225_) );
NOR2X1 NOR2X1_776 ( .A(cpuregs_11_[21]), .B(decoded_rs1_2_bF_buf5_), .Y(_9226_) );
OAI21X1 OAI21X1_1834 ( .A(_7560__bF_buf6), .B(cpuregs_15_[21]), .C(decoded_rs1_0_bF_buf52_), .Y(_9227_) );
NOR2X1 NOR2X1_777 ( .A(_9226_), .B(_9227_), .Y(_9228_) );
NOR2X1 NOR2X1_778 ( .A(cpuregs_10_[21]), .B(decoded_rs1_2_bF_buf4_), .Y(_9229_) );
OAI21X1 OAI21X1_1835 ( .A(_7560__bF_buf5), .B(cpuregs_14_[21]), .C(_7569__bF_buf9), .Y(_9230_) );
OAI21X1 OAI21X1_1836 ( .A(_9230_), .B(_9229_), .C(decoded_rs1_1_bF_buf21_), .Y(_9231_) );
NOR2X1 NOR2X1_779 ( .A(_9228_), .B(_9231_), .Y(_9232_) );
NOR2X1 NOR2X1_780 ( .A(cpuregs_9_[21]), .B(decoded_rs1_2_bF_buf3_), .Y(_9233_) );
OAI21X1 OAI21X1_1837 ( .A(_7560__bF_buf4), .B(cpuregs_13_[21]), .C(decoded_rs1_0_bF_buf51_), .Y(_9234_) );
NOR2X1 NOR2X1_781 ( .A(_9233_), .B(_9234_), .Y(_9235_) );
NOR2X1 NOR2X1_782 ( .A(cpuregs_8_[21]), .B(decoded_rs1_2_bF_buf2_), .Y(_9236_) );
OAI21X1 OAI21X1_1838 ( .A(_7560__bF_buf3), .B(cpuregs_12_[21]), .C(_7569__bF_buf8), .Y(_9237_) );
OAI21X1 OAI21X1_1839 ( .A(_9237_), .B(_9236_), .C(_7556__bF_buf21), .Y(_9238_) );
OAI21X1 OAI21X1_1840 ( .A(_9238_), .B(_9235_), .C(decoded_rs1_3_bF_buf1_), .Y(_9239_) );
INVX1 INVX1_771 ( .A(cpuregs_4_[21]), .Y(_9240_) );
OAI21X1 OAI21X1_1841 ( .A(_9240_), .B(decoded_rs1_0_bF_buf50_), .C(_7556__bF_buf20), .Y(_9241_) );
AOI21X1 AOI21X1_557 ( .A(cpuregs_5_[21]), .B(decoded_rs1_0_bF_buf49_), .C(_9241_), .Y(_9242_) );
INVX1 INVX1_772 ( .A(cpuregs_7_[21]), .Y(_9243_) );
OAI21X1 OAI21X1_1842 ( .A(_9243_), .B(_7569__bF_buf7), .C(decoded_rs1_1_bF_buf20_), .Y(_9244_) );
AOI21X1 AOI21X1_558 ( .A(cpuregs_6_[21]), .B(_7569__bF_buf6), .C(_9244_), .Y(_9245_) );
OAI21X1 OAI21X1_1843 ( .A(_9245_), .B(_9242_), .C(decoded_rs1_2_bF_buf1_), .Y(_9246_) );
INVX1 INVX1_773 ( .A(cpuregs_0_[21]), .Y(_9247_) );
OAI21X1 OAI21X1_1844 ( .A(_9247_), .B(decoded_rs1_0_bF_buf48_), .C(_7556__bF_buf19), .Y(_9248_) );
AOI21X1 AOI21X1_559 ( .A(cpuregs_1_[21]), .B(decoded_rs1_0_bF_buf47_), .C(_9248_), .Y(_9249_) );
INVX1 INVX1_774 ( .A(cpuregs_3_[21]), .Y(_9250_) );
OAI21X1 OAI21X1_1845 ( .A(_9250_), .B(_7569__bF_buf5), .C(decoded_rs1_1_bF_buf19_), .Y(_9251_) );
AOI21X1 AOI21X1_560 ( .A(cpuregs_2_[21]), .B(_7569__bF_buf4), .C(_9251_), .Y(_9252_) );
OAI21X1 OAI21X1_1846 ( .A(_9252_), .B(_9249_), .C(_7560__bF_buf2), .Y(_9253_) );
NAND3X1 NAND3X1_42 ( .A(_7561__bF_buf3), .B(_9246_), .C(_9253_), .Y(_9254_) );
OAI21X1 OAI21X1_1847 ( .A(_9232_), .B(_9239_), .C(_9254_), .Y(_9255_) );
NOR2X1 NOR2X1_783 ( .A(decoded_rs1_4_bF_buf1_), .B(_9255_), .Y(_9256_) );
NOR2X1 NOR2X1_784 ( .A(_7586__bF_buf2), .B(_9256_), .Y(_9257_) );
AOI22X1 AOI22X1_87 ( .A(reg_pc_21_), .B(_7551__bF_buf2), .C(_9257_), .D(_9225_), .Y(_9258_) );
NOR2X1 NOR2X1_785 ( .A(_4538__bF_buf3), .B(_9258_), .Y(_9259_) );
OAI21X1 OAI21X1_1848 ( .A(instr_slli), .B(instr_sll), .C(_10734__20_), .Y(_9260_) );
OAI21X1 OAI21X1_1849 ( .A(_7698__bF_buf4), .B(_9021_), .C(_9260_), .Y(_9261_) );
OAI21X1 OAI21X1_1850 ( .A(_7698__bF_buf3), .B(_5027_), .C(_9019_), .Y(_9262_) );
MUX2X1 MUX2X1_186 ( .A(_9261_), .B(_9262_), .S(_4579__bF_buf1), .Y(_9263_) );
OAI21X1 OAI21X1_1851 ( .A(_7627_), .B(_5217_), .C(resetn_bF_buf3), .Y(_9264_) );
AOI21X1 AOI21X1_561 ( .A(_10734__21_), .B(_4597__bF_buf0), .C(_9264_), .Y(_9265_) );
OAI21X1 OAI21X1_1852 ( .A(_7697__bF_buf1), .B(_9263_), .C(_9265_), .Y(_9266_) );
OR2X2 OR2X2_13 ( .A(_9259_), .B(_9266_), .Y(_9267_) );
NOR2X1 NOR2X1_786 ( .A(_9267_), .B(_9199_), .Y(_9268_) );
AOI22X1 AOI22X1_88 ( .A(_4426__bF_buf8), .B(_5217_), .C(_9268_), .D(_9197_), .Y(_81__21_) );
INVX1 INVX1_775 ( .A(decoded_imm_22_), .Y(_9269_) );
NOR2X1 NOR2X1_787 ( .A(_9021_), .B(_9269_), .Y(_9270_) );
INVX1 INVX1_776 ( .A(_9270_), .Y(_9271_) );
NAND2X1 NAND2X1_564 ( .A(_9021_), .B(_9269_), .Y(_9272_) );
NAND2X1 NAND2X1_565 ( .A(_9272_), .B(_9271_), .Y(_9273_) );
NOR2X1 NOR2X1_788 ( .A(_9110_), .B(_9191_), .Y(_9274_) );
AND2X2 AND2X2_115 ( .A(_9106_), .B(_9274_), .Y(_9275_) );
OAI21X1 OAI21X1_1853 ( .A(_9189_), .B(_9109_), .C(_9188_), .Y(_9276_) );
NOR2X1 NOR2X1_789 ( .A(_9276_), .B(_9275_), .Y(_9277_) );
NAND2X1 NAND2X1_566 ( .A(_9273_), .B(_9277_), .Y(_9278_) );
INVX1 INVX1_777 ( .A(_9273_), .Y(_9279_) );
OAI21X1 OAI21X1_1854 ( .A(_9275_), .B(_9276_), .C(_9279_), .Y(_9280_) );
NAND2X1 NAND2X1_567 ( .A(_9280_), .B(_9278_), .Y(_9281_) );
NAND2X1 NAND2X1_568 ( .A(_7624__bF_buf0), .B(_9281_), .Y(_9282_) );
AOI21X1 AOI21X1_562 ( .A(_9021_), .B(_7623__bF_buf0), .C(_4587__bF_buf0), .Y(_9283_) );
NAND2X1 NAND2X1_569 ( .A(_9283_), .B(_9282_), .Y(_9284_) );
OAI21X1 OAI21X1_1855 ( .A(_7632__bF_buf3), .B(_10734__22_), .C(_7630_), .Y(_9285_) );
AOI21X1 AOI21X1_563 ( .A(_7632__bF_buf2), .B(_9281_), .C(_9285_), .Y(_9286_) );
OAI21X1 OAI21X1_1856 ( .A(_6950_), .B(decoded_rs1_0_bF_buf46_), .C(_7556__bF_buf18), .Y(_9287_) );
AOI21X1 AOI21X1_564 ( .A(cpuregs_25_[22]), .B(decoded_rs1_0_bF_buf45_), .C(_9287_), .Y(_9288_) );
OAI21X1 OAI21X1_1857 ( .A(_6953_), .B(_7569__bF_buf3), .C(decoded_rs1_1_bF_buf18_), .Y(_9289_) );
AOI21X1 AOI21X1_565 ( .A(cpuregs_26_[22]), .B(_7569__bF_buf2), .C(_9289_), .Y(_9290_) );
OAI21X1 OAI21X1_1858 ( .A(_9288_), .B(_9290_), .C(_7560__bF_buf1), .Y(_9291_) );
OAI21X1 OAI21X1_1859 ( .A(_6942_), .B(decoded_rs1_0_bF_buf44_), .C(_7556__bF_buf17), .Y(_9292_) );
AOI21X1 AOI21X1_566 ( .A(cpuregs_29_[22]), .B(decoded_rs1_0_bF_buf43_), .C(_9292_), .Y(_9293_) );
OAI21X1 OAI21X1_1860 ( .A(_6945_), .B(_7569__bF_buf1), .C(decoded_rs1_1_bF_buf17_), .Y(_9294_) );
AOI21X1 AOI21X1_567 ( .A(cpuregs_30_[22]), .B(_7569__bF_buf0), .C(_9294_), .Y(_9295_) );
OAI21X1 OAI21X1_1861 ( .A(_9293_), .B(_9295_), .C(decoded_rs1_2_bF_buf0_), .Y(_9296_) );
AOI21X1 AOI21X1_568 ( .A(_9291_), .B(_9296_), .C(_7561__bF_buf2), .Y(_9297_) );
MUX2X1 MUX2X1_187 ( .A(cpuregs_22_[22]), .B(cpuregs_20_[22]), .S(decoded_rs1_1_bF_buf16_), .Y(_9298_) );
NAND2X1 NAND2X1_570 ( .A(cpuregs_23_[22]), .B(decoded_rs1_1_bF_buf15_), .Y(_9299_) );
OAI21X1 OAI21X1_1862 ( .A(_6965_), .B(decoded_rs1_1_bF_buf14_), .C(_9299_), .Y(_9300_) );
AOI21X1 AOI21X1_569 ( .A(decoded_rs1_0_bF_buf42_), .B(_9300_), .C(_7560__bF_buf0), .Y(_9301_) );
OAI21X1 OAI21X1_1863 ( .A(decoded_rs1_0_bF_buf41_), .B(_9298_), .C(_9301_), .Y(_9302_) );
MUX2X1 MUX2X1_188 ( .A(cpuregs_18_[22]), .B(cpuregs_16_[22]), .S(decoded_rs1_1_bF_buf13_), .Y(_9303_) );
NAND2X1 NAND2X1_571 ( .A(cpuregs_19_[22]), .B(decoded_rs1_1_bF_buf12_), .Y(_9304_) );
OAI21X1 OAI21X1_1864 ( .A(_6959_), .B(decoded_rs1_1_bF_buf11_), .C(_9304_), .Y(_9305_) );
AOI21X1 AOI21X1_570 ( .A(decoded_rs1_0_bF_buf40_), .B(_9305_), .C(decoded_rs1_2_bF_buf12_), .Y(_9306_) );
OAI21X1 OAI21X1_1865 ( .A(decoded_rs1_0_bF_buf39_), .B(_9303_), .C(_9306_), .Y(_9307_) );
AOI21X1 AOI21X1_571 ( .A(_9302_), .B(_9307_), .C(decoded_rs1_3_bF_buf0_), .Y(_9308_) );
OAI21X1 OAI21X1_1866 ( .A(_9297_), .B(_9308_), .C(decoded_rs1_4_bF_buf0_), .Y(_9309_) );
AOI21X1 AOI21X1_572 ( .A(_6934_), .B(_7556__bF_buf16), .C(_7569__bF_buf48), .Y(_9310_) );
OAI21X1 OAI21X1_1867 ( .A(cpuregs_15_[22]), .B(_7556__bF_buf15), .C(_9310_), .Y(_9311_) );
INVX1 INVX1_778 ( .A(cpuregs_12_[22]), .Y(_9312_) );
AOI21X1 AOI21X1_573 ( .A(_9312_), .B(_7556__bF_buf14), .C(decoded_rs1_0_bF_buf38_), .Y(_9313_) );
OAI21X1 OAI21X1_1868 ( .A(cpuregs_14_[22]), .B(_7556__bF_buf13), .C(_9313_), .Y(_9314_) );
NAND3X1 NAND3X1_43 ( .A(decoded_rs1_2_bF_buf11_), .B(_9311_), .C(_9314_), .Y(_9315_) );
AND2X2 AND2X2_116 ( .A(cpuregs_9_[22]), .B(decoded_rs1_0_bF_buf37_), .Y(_9316_) );
INVX1 INVX1_779 ( .A(cpuregs_8_[22]), .Y(_9317_) );
OAI21X1 OAI21X1_1869 ( .A(_9317_), .B(decoded_rs1_0_bF_buf36_), .C(_7556__bF_buf12), .Y(_9318_) );
INVX1 INVX1_780 ( .A(cpuregs_10_[22]), .Y(_9319_) );
AOI21X1 AOI21X1_574 ( .A(cpuregs_11_[22]), .B(decoded_rs1_0_bF_buf35_), .C(_7556__bF_buf11), .Y(_9320_) );
OAI21X1 OAI21X1_1870 ( .A(_9319_), .B(decoded_rs1_0_bF_buf34_), .C(_9320_), .Y(_9321_) );
OAI21X1 OAI21X1_1871 ( .A(_9316_), .B(_9318_), .C(_9321_), .Y(_9322_) );
AOI21X1 AOI21X1_575 ( .A(_7560__bF_buf12), .B(_9322_), .C(_7561__bF_buf1), .Y(_9323_) );
INVX1 INVX1_781 ( .A(cpuregs_7_[22]), .Y(_9324_) );
AOI21X1 AOI21X1_576 ( .A(decoded_rs1_2_bF_buf10_), .B(_9324_), .C(_7569__bF_buf47), .Y(_9325_) );
OAI21X1 OAI21X1_1872 ( .A(cpuregs_3_[22]), .B(decoded_rs1_2_bF_buf9_), .C(_9325_), .Y(_9326_) );
OAI21X1 OAI21X1_1873 ( .A(_7560__bF_buf11), .B(cpuregs_6_[22]), .C(_7569__bF_buf46), .Y(_9327_) );
AOI21X1 AOI21X1_577 ( .A(_6922_), .B(_7560__bF_buf10), .C(_9327_), .Y(_9328_) );
NOR2X1 NOR2X1_790 ( .A(_7556__bF_buf10), .B(_9328_), .Y(_9329_) );
NOR2X1 NOR2X1_791 ( .A(cpuregs_1_[22]), .B(decoded_rs1_2_bF_buf8_), .Y(_9330_) );
OAI21X1 OAI21X1_1874 ( .A(_7560__bF_buf9), .B(cpuregs_5_[22]), .C(decoded_rs1_0_bF_buf33_), .Y(_9331_) );
NOR2X1 NOR2X1_792 ( .A(_9330_), .B(_9331_), .Y(_9332_) );
NOR2X1 NOR2X1_793 ( .A(cpuregs_0_[22]), .B(decoded_rs1_2_bF_buf7_), .Y(_9333_) );
OAI21X1 OAI21X1_1875 ( .A(_7560__bF_buf8), .B(cpuregs_4_[22]), .C(_7569__bF_buf45), .Y(_9334_) );
OAI21X1 OAI21X1_1876 ( .A(_9334_), .B(_9333_), .C(_7556__bF_buf9), .Y(_9335_) );
OAI21X1 OAI21X1_1877 ( .A(_9335_), .B(_9332_), .C(_7561__bF_buf0), .Y(_9336_) );
AOI21X1 AOI21X1_578 ( .A(_9326_), .B(_9329_), .C(_9336_), .Y(_9337_) );
AOI21X1 AOI21X1_579 ( .A(_9315_), .B(_9323_), .C(_9337_), .Y(_9338_) );
AOI21X1 AOI21X1_580 ( .A(_7552__bF_buf1), .B(_9338_), .C(_7586__bF_buf1), .Y(_9339_) );
AOI22X1 AOI22X1_89 ( .A(reg_pc_22_), .B(_7551__bF_buf1), .C(_9339_), .D(_9309_), .Y(_9340_) );
NOR2X1 NOR2X1_794 ( .A(_4538__bF_buf2), .B(_9340_), .Y(_9341_) );
NOR2X1 NOR2X1_795 ( .A(_5045_), .B(_7700__bF_buf5), .Y(_9342_) );
OAI21X1 OAI21X1_1878 ( .A(instr_slli), .B(instr_sll), .C(_10734__21_), .Y(_9343_) );
OAI21X1 OAI21X1_1879 ( .A(_7698__bF_buf2), .B(_9091_), .C(_9343_), .Y(_9344_) );
OAI21X1 OAI21X1_1880 ( .A(_7698__bF_buf1), .B(_5021_), .C(_4580__bF_buf2), .Y(_9345_) );
OAI22X1 OAI22X1_186 ( .A(_4580__bF_buf1), .B(_9344_), .C(_9345_), .D(_9342_), .Y(_9346_) );
OAI21X1 OAI21X1_1881 ( .A(_7627_), .B(_9021_), .C(resetn_bF_buf2), .Y(_9347_) );
AOI21X1 AOI21X1_581 ( .A(_10734__22_), .B(_4597__bF_buf3), .C(_9347_), .Y(_9348_) );
OAI21X1 OAI21X1_1882 ( .A(_7697__bF_buf0), .B(_9346_), .C(_9348_), .Y(_9349_) );
OR2X2 OR2X2_14 ( .A(_9341_), .B(_9349_), .Y(_9350_) );
NOR2X1 NOR2X1_796 ( .A(_9350_), .B(_9286_), .Y(_9351_) );
AOI22X1 AOI22X1_90 ( .A(_4426__bF_buf7), .B(_9021_), .C(_9351_), .D(_9284_), .Y(_81__22_) );
NAND2X1 NAND2X1_572 ( .A(_10734__23_), .B(decoded_imm_23_), .Y(_9352_) );
NOR2X1 NOR2X1_797 ( .A(_10734__23_), .B(decoded_imm_23_), .Y(_9353_) );
INVX1 INVX1_782 ( .A(_9353_), .Y(_9354_) );
NAND2X1 NAND2X1_573 ( .A(_9352_), .B(_9354_), .Y(_9355_) );
INVX1 INVX1_783 ( .A(_9355_), .Y(_9356_) );
NAND3X1 NAND3X1_44 ( .A(_9271_), .B(_9356_), .C(_9280_), .Y(_9357_) );
OAI21X1 OAI21X1_1883 ( .A(_9021_), .B(_9269_), .C(_9280_), .Y(_9358_) );
INVX1 INVX1_784 ( .A(_9352_), .Y(_9359_) );
OAI21X1 OAI21X1_1884 ( .A(_9359_), .B(_9353_), .C(_9358_), .Y(_9360_) );
NAND2X1 NAND2X1_574 ( .A(_9357_), .B(_9360_), .Y(_9361_) );
AOI21X1 AOI21X1_582 ( .A(_9091_), .B(_7623__bF_buf4), .C(_4587__bF_buf3), .Y(_9362_) );
OAI21X1 OAI21X1_1885 ( .A(_9361_), .B(_7623__bF_buf3), .C(_9362_), .Y(_9363_) );
NAND3X1 NAND3X1_45 ( .A(_7632__bF_buf1), .B(_9357_), .C(_9360_), .Y(_9364_) );
AOI21X1 AOI21X1_583 ( .A(_9091_), .B(_7631__bF_buf3), .C(_7629__bF_buf0), .Y(_9365_) );
OAI21X1 OAI21X1_1886 ( .A(_7007_), .B(decoded_rs1_0_bF_buf32_), .C(_7556__bF_buf8), .Y(_9366_) );
AOI21X1 AOI21X1_584 ( .A(cpuregs_17_[23]), .B(decoded_rs1_0_bF_buf31_), .C(_9366_), .Y(_9367_) );
NAND2X1 NAND2X1_575 ( .A(_7010_), .B(_7569__bF_buf44), .Y(_9368_) );
OAI21X1 OAI21X1_1887 ( .A(cpuregs_19_[23]), .B(_7569__bF_buf43), .C(_9368_), .Y(_9369_) );
AOI21X1 AOI21X1_585 ( .A(decoded_rs1_1_bF_buf10_), .B(_9369_), .C(_9367_), .Y(_9370_) );
AND2X2 AND2X2_117 ( .A(cpuregs_21_[23]), .B(decoded_rs1_0_bF_buf30_), .Y(_9371_) );
OAI21X1 OAI21X1_1888 ( .A(_7014_), .B(decoded_rs1_0_bF_buf29_), .C(_7556__bF_buf7), .Y(_9372_) );
AOI21X1 AOI21X1_586 ( .A(cpuregs_23_[23]), .B(decoded_rs1_0_bF_buf28_), .C(_7556__bF_buf6), .Y(_9373_) );
OAI21X1 OAI21X1_1889 ( .A(_7017_), .B(decoded_rs1_0_bF_buf27_), .C(_9373_), .Y(_9374_) );
OAI21X1 OAI21X1_1890 ( .A(_9371_), .B(_9372_), .C(_9374_), .Y(_9375_) );
OAI21X1 OAI21X1_1891 ( .A(_9375_), .B(_7560__bF_buf7), .C(_7561__bF_buf6), .Y(_9376_) );
AOI21X1 AOI21X1_587 ( .A(_7560__bF_buf6), .B(_9370_), .C(_9376_), .Y(_9377_) );
OAI21X1 OAI21X1_1892 ( .A(cpuregs_25_[23]), .B(decoded_rs1_1_bF_buf9_), .C(decoded_rs1_0_bF_buf26_), .Y(_9378_) );
AOI21X1 AOI21X1_588 ( .A(_7033_), .B(decoded_rs1_1_bF_buf8_), .C(_9378_), .Y(_9379_) );
NOR2X1 NOR2X1_798 ( .A(cpuregs_26_[23]), .B(_7556__bF_buf5), .Y(_9380_) );
OAI21X1 OAI21X1_1893 ( .A(cpuregs_24_[23]), .B(decoded_rs1_1_bF_buf7_), .C(_7569__bF_buf42), .Y(_9381_) );
OAI21X1 OAI21X1_1894 ( .A(_9380_), .B(_9381_), .C(_7560__bF_buf5), .Y(_9382_) );
OAI21X1 OAI21X1_1895 ( .A(cpuregs_29_[23]), .B(decoded_rs1_1_bF_buf6_), .C(decoded_rs1_0_bF_buf25_), .Y(_9383_) );
AOI21X1 AOI21X1_589 ( .A(_7025_), .B(decoded_rs1_1_bF_buf5_), .C(_9383_), .Y(_9384_) );
NOR2X1 NOR2X1_799 ( .A(cpuregs_30_[23]), .B(_7556__bF_buf4), .Y(_9385_) );
OAI21X1 OAI21X1_1896 ( .A(cpuregs_28_[23]), .B(decoded_rs1_1_bF_buf4_), .C(_7569__bF_buf41), .Y(_9386_) );
OAI21X1 OAI21X1_1897 ( .A(_9385_), .B(_9386_), .C(decoded_rs1_2_bF_buf6_), .Y(_9387_) );
OAI22X1 OAI22X1_187 ( .A(_9382_), .B(_9379_), .C(_9384_), .D(_9387_), .Y(_9388_) );
AND2X2 AND2X2_118 ( .A(_9388_), .B(decoded_rs1_3_bF_buf6_), .Y(_9389_) );
OAI21X1 OAI21X1_1898 ( .A(_9377_), .B(_9389_), .C(decoded_rs1_4_bF_buf4_), .Y(_9390_) );
AND2X2 AND2X2_119 ( .A(cpuregs_9_[23]), .B(decoded_rs1_0_bF_buf24_), .Y(_9391_) );
OAI21X1 OAI21X1_1899 ( .A(_6991_), .B(decoded_rs1_0_bF_buf23_), .C(_7556__bF_buf3), .Y(_9392_) );
AOI21X1 AOI21X1_590 ( .A(cpuregs_11_[23]), .B(decoded_rs1_0_bF_buf22_), .C(_7556__bF_buf2), .Y(_9393_) );
OAI21X1 OAI21X1_1900 ( .A(_6994_), .B(decoded_rs1_0_bF_buf21_), .C(_9393_), .Y(_9394_) );
OAI21X1 OAI21X1_1901 ( .A(_9391_), .B(_9392_), .C(_9394_), .Y(_9395_) );
AOI21X1 AOI21X1_591 ( .A(cpuregs_12_[23]), .B(_7569__bF_buf40), .C(decoded_rs1_1_bF_buf3_), .Y(_9396_) );
OAI21X1 OAI21X1_1902 ( .A(_6999_), .B(_7569__bF_buf39), .C(_9396_), .Y(_9397_) );
INVX1 INVX1_785 ( .A(cpuregs_14_[23]), .Y(_9398_) );
AOI21X1 AOI21X1_592 ( .A(cpuregs_15_[23]), .B(decoded_rs1_0_bF_buf20_), .C(_7556__bF_buf1), .Y(_9399_) );
OAI21X1 OAI21X1_1903 ( .A(_9398_), .B(decoded_rs1_0_bF_buf19_), .C(_9399_), .Y(_9400_) );
AOI21X1 AOI21X1_593 ( .A(_9397_), .B(_9400_), .C(_7560__bF_buf4), .Y(_9401_) );
AOI21X1 AOI21X1_594 ( .A(_7560__bF_buf3), .B(_9395_), .C(_9401_), .Y(_9402_) );
AND2X2 AND2X2_120 ( .A(cpuregs_5_[23]), .B(decoded_rs1_0_bF_buf18_), .Y(_9403_) );
INVX1 INVX1_786 ( .A(cpuregs_4_[23]), .Y(_9404_) );
OAI21X1 OAI21X1_1904 ( .A(_9404_), .B(decoded_rs1_0_bF_buf17_), .C(_7556__bF_buf0), .Y(_9405_) );
NOR2X1 NOR2X1_800 ( .A(decoded_rs1_0_bF_buf16_), .B(_6986_), .Y(_9406_) );
INVX1 INVX1_787 ( .A(cpuregs_7_[23]), .Y(_9407_) );
OAI21X1 OAI21X1_1905 ( .A(_9407_), .B(_7569__bF_buf38), .C(decoded_rs1_1_bF_buf2_), .Y(_9408_) );
OAI22X1 OAI22X1_188 ( .A(_9405_), .B(_9403_), .C(_9408_), .D(_9406_), .Y(_9409_) );
AOI21X1 AOI21X1_595 ( .A(cpuregs_0_[23]), .B(_7569__bF_buf37), .C(decoded_rs1_1_bF_buf1_), .Y(_9410_) );
OAI21X1 OAI21X1_1906 ( .A(_6978_), .B(_7569__bF_buf36), .C(_9410_), .Y(_9411_) );
INVX1 INVX1_788 ( .A(cpuregs_2_[23]), .Y(_9412_) );
AOI21X1 AOI21X1_596 ( .A(cpuregs_3_[23]), .B(decoded_rs1_0_bF_buf15_), .C(_7556__bF_buf42), .Y(_9413_) );
OAI21X1 OAI21X1_1907 ( .A(_9412_), .B(decoded_rs1_0_bF_buf14_), .C(_9413_), .Y(_9414_) );
NAND3X1 NAND3X1_46 ( .A(_7560__bF_buf2), .B(_9411_), .C(_9414_), .Y(_9415_) );
OAI21X1 OAI21X1_1908 ( .A(_7560__bF_buf1), .B(_9409_), .C(_9415_), .Y(_9416_) );
MUX2X1 MUX2X1_189 ( .A(_9402_), .B(_9416_), .S(decoded_rs1_3_bF_buf5_), .Y(_9417_) );
AOI21X1 AOI21X1_597 ( .A(_7552__bF_buf0), .B(_9417_), .C(_7586__bF_buf0), .Y(_9418_) );
AOI22X1 AOI22X1_91 ( .A(reg_pc_23_), .B(_7551__bF_buf0), .C(_9418_), .D(_9390_), .Y(_9419_) );
OAI21X1 OAI21X1_1909 ( .A(instr_slli), .B(instr_sll), .C(_10734__22_), .Y(_9420_) );
OAI21X1 OAI21X1_1910 ( .A(_7698__bF_buf0), .B(_5032_), .C(_9420_), .Y(_9421_) );
NAND2X1 NAND2X1_576 ( .A(_4579__bF_buf0), .B(_9421_), .Y(_9422_) );
NOR2X1 NOR2X1_801 ( .A(_5016_), .B(_7698__bF_buf4), .Y(_9423_) );
OAI21X1 OAI21X1_1911 ( .A(_9423_), .B(_9183_), .C(_4580__bF_buf0), .Y(_9424_) );
NAND2X1 NAND2X1_577 ( .A(_9422_), .B(_9424_), .Y(_9425_) );
NAND2X1 NAND2X1_578 ( .A(_9425_), .B(_4584_), .Y(_9426_) );
OAI21X1 OAI21X1_1912 ( .A(_7627_), .B(_9091_), .C(resetn_bF_buf1), .Y(_9427_) );
AOI21X1 AOI21X1_598 ( .A(_10734__23_), .B(_4597__bF_buf2), .C(_9427_), .Y(_9428_) );
AND2X2 AND2X2_121 ( .A(_9426_), .B(_9428_), .Y(_9429_) );
OAI21X1 OAI21X1_1913 ( .A(_9419_), .B(_4538__bF_buf1), .C(_9429_), .Y(_9430_) );
AOI21X1 AOI21X1_599 ( .A(_9365_), .B(_9364_), .C(_9430_), .Y(_9431_) );
AOI22X1 AOI22X1_92 ( .A(_4426__bF_buf6), .B(_9091_), .C(_9431_), .D(_9363_), .Y(_81__23_) );
NOR2X1 NOR2X1_802 ( .A(_9355_), .B(_9273_), .Y(_9432_) );
NAND2X1 NAND2X1_579 ( .A(_9274_), .B(_9432_), .Y(_9433_) );
OAI21X1 OAI21X1_1914 ( .A(_9270_), .B(_9359_), .C(_9354_), .Y(_9434_) );
OAI21X1 OAI21X1_1915 ( .A(_9103_), .B(_9433_), .C(_9434_), .Y(_9435_) );
AOI21X1 AOI21X1_600 ( .A(_9276_), .B(_9432_), .C(_9435_), .Y(_9436_) );
NOR2X1 NOR2X1_803 ( .A(_9433_), .B(_9105_), .Y(_9437_) );
INVX1 INVX1_789 ( .A(_9437_), .Y(_9438_) );
OAI21X1 OAI21X1_1916 ( .A(_8781_), .B(_9438_), .C(_9436_), .Y(_9439_) );
INVX1 INVX1_790 ( .A(decoded_imm_24_), .Y(_9440_) );
NAND2X1 NAND2X1_580 ( .A(_5032_), .B(_9440_), .Y(_9441_) );
NOR2X1 NOR2X1_804 ( .A(_5032_), .B(_9440_), .Y(_9442_) );
INVX1 INVX1_791 ( .A(_9442_), .Y(_9443_) );
AND2X2 AND2X2_122 ( .A(_9443_), .B(_9441_), .Y(_9444_) );
XNOR2X1 XNOR2X1_13 ( .A(_9439_), .B(_9444_), .Y(_9445_) );
OAI21X1 OAI21X1_1917 ( .A(_7632__bF_buf0), .B(_10734__24_), .C(_7630_), .Y(_9446_) );
AOI21X1 AOI21X1_601 ( .A(_7632__bF_buf3), .B(_9445_), .C(_9446_), .Y(_9447_) );
INVX1 INVX1_792 ( .A(_9445_), .Y(_9448_) );
NOR2X1 NOR2X1_805 ( .A(_7623__bF_buf2), .B(_9448_), .Y(_9449_) );
OAI21X1 OAI21X1_1918 ( .A(_7624__bF_buf4), .B(_10734__24_), .C(cpu_state_5_bF_buf2_), .Y(_9450_) );
OAI21X1 OAI21X1_1919 ( .A(_7070_), .B(decoded_rs1_0_bF_buf13_), .C(_7556__bF_buf41), .Y(_9451_) );
AOI21X1 AOI21X1_602 ( .A(cpuregs_17_[24]), .B(decoded_rs1_0_bF_buf12_), .C(_9451_), .Y(_9452_) );
NAND2X1 NAND2X1_581 ( .A(_7073_), .B(_7569__bF_buf35), .Y(_9453_) );
OAI21X1 OAI21X1_1920 ( .A(cpuregs_19_[24]), .B(_7569__bF_buf34), .C(_9453_), .Y(_9454_) );
AOI21X1 AOI21X1_603 ( .A(decoded_rs1_1_bF_buf0_), .B(_9454_), .C(_9452_), .Y(_9455_) );
AND2X2 AND2X2_123 ( .A(cpuregs_21_[24]), .B(decoded_rs1_0_bF_buf11_), .Y(_9456_) );
OAI21X1 OAI21X1_1921 ( .A(_7077_), .B(decoded_rs1_0_bF_buf10_), .C(_7556__bF_buf40), .Y(_9457_) );
AOI21X1 AOI21X1_604 ( .A(cpuregs_23_[24]), .B(decoded_rs1_0_bF_buf9_), .C(_7556__bF_buf39), .Y(_9458_) );
OAI21X1 OAI21X1_1922 ( .A(_7080_), .B(decoded_rs1_0_bF_buf8_), .C(_9458_), .Y(_9459_) );
OAI21X1 OAI21X1_1923 ( .A(_9456_), .B(_9457_), .C(_9459_), .Y(_9460_) );
OAI21X1 OAI21X1_1924 ( .A(_9460_), .B(_7560__bF_buf0), .C(_7561__bF_buf5), .Y(_9461_) );
AOI21X1 AOI21X1_605 ( .A(_7560__bF_buf12), .B(_9455_), .C(_9461_), .Y(_9462_) );
OAI21X1 OAI21X1_1925 ( .A(cpuregs_25_[24]), .B(decoded_rs1_1_bF_buf44_), .C(decoded_rs1_0_bF_buf7_), .Y(_9463_) );
AOI21X1 AOI21X1_606 ( .A(_7096_), .B(decoded_rs1_1_bF_buf43_), .C(_9463_), .Y(_9464_) );
NOR2X1 NOR2X1_806 ( .A(cpuregs_26_[24]), .B(_7556__bF_buf38), .Y(_9465_) );
OAI21X1 OAI21X1_1926 ( .A(cpuregs_24_[24]), .B(decoded_rs1_1_bF_buf42_), .C(_7569__bF_buf33), .Y(_9466_) );
OAI21X1 OAI21X1_1927 ( .A(_9465_), .B(_9466_), .C(_7560__bF_buf11), .Y(_9467_) );
OAI21X1 OAI21X1_1928 ( .A(cpuregs_29_[24]), .B(decoded_rs1_1_bF_buf41_), .C(decoded_rs1_0_bF_buf6_), .Y(_9468_) );
AOI21X1 AOI21X1_607 ( .A(_7088_), .B(decoded_rs1_1_bF_buf40_), .C(_9468_), .Y(_9469_) );
NOR2X1 NOR2X1_807 ( .A(cpuregs_30_[24]), .B(_7556__bF_buf37), .Y(_9470_) );
OAI21X1 OAI21X1_1929 ( .A(cpuregs_28_[24]), .B(decoded_rs1_1_bF_buf39_), .C(_7569__bF_buf32), .Y(_9471_) );
OAI21X1 OAI21X1_1930 ( .A(_9470_), .B(_9471_), .C(decoded_rs1_2_bF_buf5_), .Y(_9472_) );
OAI22X1 OAI22X1_189 ( .A(_9467_), .B(_9464_), .C(_9469_), .D(_9472_), .Y(_9473_) );
AND2X2 AND2X2_124 ( .A(_9473_), .B(decoded_rs1_3_bF_buf4_), .Y(_9474_) );
OAI21X1 OAI21X1_1931 ( .A(_9462_), .B(_9474_), .C(decoded_rs1_4_bF_buf3_), .Y(_9475_) );
AND2X2 AND2X2_125 ( .A(cpuregs_5_[24]), .B(decoded_rs1_0_bF_buf5_), .Y(_9476_) );
INVX1 INVX1_793 ( .A(cpuregs_4_[24]), .Y(_9477_) );
OAI21X1 OAI21X1_1932 ( .A(_9477_), .B(decoded_rs1_0_bF_buf4_), .C(_7556__bF_buf36), .Y(_9478_) );
NOR2X1 NOR2X1_808 ( .A(decoded_rs1_0_bF_buf3_), .B(_7049_), .Y(_9479_) );
INVX1 INVX1_794 ( .A(cpuregs_7_[24]), .Y(_9480_) );
OAI21X1 OAI21X1_1933 ( .A(_9480_), .B(_7569__bF_buf31), .C(decoded_rs1_1_bF_buf38_), .Y(_9481_) );
OAI22X1 OAI22X1_190 ( .A(_9478_), .B(_9476_), .C(_9481_), .D(_9479_), .Y(_9482_) );
AOI21X1 AOI21X1_608 ( .A(cpuregs_0_[24]), .B(_7569__bF_buf30), .C(decoded_rs1_1_bF_buf37_), .Y(_9483_) );
OAI21X1 OAI21X1_1934 ( .A(_7042_), .B(_7569__bF_buf29), .C(_9483_), .Y(_9484_) );
INVX1 INVX1_795 ( .A(cpuregs_2_[24]), .Y(_9485_) );
AOI21X1 AOI21X1_609 ( .A(cpuregs_3_[24]), .B(decoded_rs1_0_bF_buf2_), .C(_7556__bF_buf35), .Y(_9486_) );
OAI21X1 OAI21X1_1935 ( .A(_9485_), .B(decoded_rs1_0_bF_buf1_), .C(_9486_), .Y(_9487_) );
NAND3X1 NAND3X1_47 ( .A(_7560__bF_buf10), .B(_9484_), .C(_9487_), .Y(_9488_) );
OAI21X1 OAI21X1_1936 ( .A(_7560__bF_buf9), .B(_9482_), .C(_9488_), .Y(_9489_) );
OAI21X1 OAI21X1_1937 ( .A(_7560__bF_buf8), .B(cpuregs_13_[24]), .C(decoded_rs1_0_bF_buf0_), .Y(_9490_) );
AOI21X1 AOI21X1_610 ( .A(_7062_), .B(_7560__bF_buf7), .C(_9490_), .Y(_9491_) );
NOR2X1 NOR2X1_809 ( .A(cpuregs_8_[24]), .B(decoded_rs1_2_bF_buf4_), .Y(_9492_) );
OAI21X1 OAI21X1_1938 ( .A(_7560__bF_buf6), .B(cpuregs_12_[24]), .C(_7569__bF_buf28), .Y(_9493_) );
OAI21X1 OAI21X1_1939 ( .A(_9493_), .B(_9492_), .C(_7556__bF_buf34), .Y(_9494_) );
NOR2X1 NOR2X1_810 ( .A(_9491_), .B(_9494_), .Y(_9495_) );
NOR2X1 NOR2X1_811 ( .A(cpuregs_11_[24]), .B(decoded_rs1_2_bF_buf3_), .Y(_9496_) );
OAI21X1 OAI21X1_1940 ( .A(_7560__bF_buf5), .B(cpuregs_15_[24]), .C(decoded_rs1_0_bF_buf57_), .Y(_9497_) );
NOR2X1 NOR2X1_812 ( .A(_9496_), .B(_9497_), .Y(_9498_) );
NOR2X1 NOR2X1_813 ( .A(cpuregs_10_[24]), .B(decoded_rs1_2_bF_buf2_), .Y(_9499_) );
OAI21X1 OAI21X1_1941 ( .A(_7560__bF_buf4), .B(cpuregs_14_[24]), .C(_7569__bF_buf27), .Y(_9500_) );
OAI21X1 OAI21X1_1942 ( .A(_9500_), .B(_9499_), .C(decoded_rs1_1_bF_buf36_), .Y(_9501_) );
NOR2X1 NOR2X1_814 ( .A(_9498_), .B(_9501_), .Y(_9502_) );
OAI21X1 OAI21X1_1943 ( .A(_9495_), .B(_9502_), .C(decoded_rs1_3_bF_buf3_), .Y(_9503_) );
OAI21X1 OAI21X1_1944 ( .A(decoded_rs1_3_bF_buf2_), .B(_9489_), .C(_9503_), .Y(_9504_) );
AOI21X1 AOI21X1_611 ( .A(_7552__bF_buf5), .B(_9504_), .C(_7586__bF_buf3), .Y(_9505_) );
NAND2X1 NAND2X1_582 ( .A(_9475_), .B(_9505_), .Y(_9506_) );
OAI21X1 OAI21X1_1945 ( .A(_4841_), .B(_7643_), .C(_9506_), .Y(_9507_) );
OAI21X1 OAI21X1_1946 ( .A(_7698__bF_buf3), .B(_5004_), .C(_9260_), .Y(_9508_) );
NOR2X1 NOR2X1_815 ( .A(_4579__bF_buf4), .B(_9508_), .Y(_9509_) );
OAI21X1 OAI21X1_1947 ( .A(instr_slli), .B(instr_sll), .C(_10734__23_), .Y(_9510_) );
OAI21X1 OAI21X1_1948 ( .A(_7698__bF_buf2), .B(_5027_), .C(_9510_), .Y(_9511_) );
NOR2X1 NOR2X1_816 ( .A(_4580__bF_buf4), .B(_9511_), .Y(_9512_) );
OAI21X1 OAI21X1_1949 ( .A(_9509_), .B(_9512_), .C(_4582_), .Y(_9513_) );
OAI21X1 OAI21X1_1950 ( .A(_10734__24_), .B(_4582_), .C(_9513_), .Y(_9514_) );
OAI22X1 OAI22X1_191 ( .A(_5032_), .B(_7627_), .C(_9514_), .D(_4575__bF_buf2), .Y(_9515_) );
AOI21X1 AOI21X1_612 ( .A(cpu_state_2_bF_buf5_), .B(_9507_), .C(_9515_), .Y(_9516_) );
OAI21X1 OAI21X1_1951 ( .A(_9449_), .B(_9450_), .C(_9516_), .Y(_9517_) );
OAI21X1 OAI21X1_1952 ( .A(_9517_), .B(_9447_), .C(resetn_bF_buf0), .Y(_9518_) );
OAI21X1 OAI21X1_1953 ( .A(resetn_bF_buf11), .B(_5032_), .C(_9518_), .Y(_81__24_) );
NOR2X1 NOR2X1_817 ( .A(_10734__25_), .B(decoded_imm_25_), .Y(_9519_) );
INVX1 INVX1_796 ( .A(decoded_imm_25_), .Y(_9520_) );
NOR2X1 NOR2X1_818 ( .A(_5027_), .B(_9520_), .Y(_9521_) );
OAI21X1 OAI21X1_1954 ( .A(_9519_), .B(_9521_), .C(_9443_), .Y(_9522_) );
AOI21X1 AOI21X1_613 ( .A(_9444_), .B(_9439_), .C(_9522_), .Y(_9523_) );
NOR2X1 NOR2X1_819 ( .A(_9519_), .B(_9521_), .Y(_9524_) );
INVX1 INVX1_797 ( .A(_9524_), .Y(_9525_) );
NOR2X1 NOR2X1_820 ( .A(_9443_), .B(_9525_), .Y(_9526_) );
NAND2X1 NAND2X1_583 ( .A(_8779_), .B(_8780_), .Y(_9527_) );
NAND2X1 NAND2X1_584 ( .A(_9437_), .B(_9527_), .Y(_9528_) );
AND2X2 AND2X2_126 ( .A(_9444_), .B(_9524_), .Y(_9529_) );
INVX1 INVX1_798 ( .A(_9529_), .Y(_9530_) );
AOI21X1 AOI21X1_614 ( .A(_9436_), .B(_9528_), .C(_9530_), .Y(_9531_) );
OR2X2 OR2X2_15 ( .A(_9531_), .B(_9526_), .Y(_9532_) );
OAI21X1 OAI21X1_1955 ( .A(_9532_), .B(_9523_), .C(_7632__bF_buf2), .Y(_9533_) );
AOI21X1 AOI21X1_615 ( .A(_5027_), .B(_7631__bF_buf2), .C(_7629__bF_buf3), .Y(_9534_) );
NAND2X1 NAND2X1_585 ( .A(_9534_), .B(_9533_), .Y(_9535_) );
OAI21X1 OAI21X1_1956 ( .A(_9532_), .B(_9523_), .C(_7624__bF_buf3), .Y(_9536_) );
AOI21X1 AOI21X1_616 ( .A(_5027_), .B(_7623__bF_buf1), .C(_4587__bF_buf2), .Y(_9537_) );
AOI21X1 AOI21X1_617 ( .A(decoded_rs1_2_bF_buf1_), .B(_7142_), .C(_7569__bF_buf26), .Y(_9538_) );
OAI21X1 OAI21X1_1957 ( .A(cpuregs_25_[25]), .B(decoded_rs1_2_bF_buf0_), .C(_9538_), .Y(_9539_) );
OAI21X1 OAI21X1_1958 ( .A(_7560__bF_buf3), .B(cpuregs_28_[25]), .C(_7569__bF_buf25), .Y(_9540_) );
AOI21X1 AOI21X1_618 ( .A(_7139_), .B(_7560__bF_buf2), .C(_9540_), .Y(_9541_) );
NOR2X1 NOR2X1_821 ( .A(decoded_rs1_1_bF_buf35_), .B(_9541_), .Y(_9542_) );
AOI21X1 AOI21X1_619 ( .A(decoded_rs1_2_bF_buf12_), .B(_7145_), .C(_7569__bF_buf24), .Y(_9543_) );
OAI21X1 OAI21X1_1959 ( .A(cpuregs_27_[25]), .B(decoded_rs1_2_bF_buf11_), .C(_9543_), .Y(_9544_) );
OAI21X1 OAI21X1_1960 ( .A(_7560__bF_buf1), .B(cpuregs_30_[25]), .C(_7569__bF_buf23), .Y(_9545_) );
AOI21X1 AOI21X1_620 ( .A(_7135_), .B(_7560__bF_buf0), .C(_9545_), .Y(_9546_) );
NOR2X1 NOR2X1_822 ( .A(_7556__bF_buf33), .B(_9546_), .Y(_9547_) );
AOI22X1 AOI22X1_93 ( .A(_9542_), .B(_9539_), .C(_9544_), .D(_9547_), .Y(_9548_) );
INVX1 INVX1_799 ( .A(cpuregs_11_[25]), .Y(_9549_) );
OAI21X1 OAI21X1_1961 ( .A(cpuregs_9_[25]), .B(decoded_rs1_1_bF_buf34_), .C(decoded_rs1_0_bF_buf56_), .Y(_9550_) );
AOI21X1 AOI21X1_621 ( .A(_9549_), .B(decoded_rs1_1_bF_buf33_), .C(_9550_), .Y(_9551_) );
NOR2X1 NOR2X1_823 ( .A(cpuregs_10_[25]), .B(_7556__bF_buf32), .Y(_9552_) );
OAI21X1 OAI21X1_1962 ( .A(cpuregs_8_[25]), .B(decoded_rs1_1_bF_buf32_), .C(_7569__bF_buf22), .Y(_9553_) );
OAI21X1 OAI21X1_1963 ( .A(_9552_), .B(_9553_), .C(_7560__bF_buf12), .Y(_9554_) );
OAI21X1 OAI21X1_1964 ( .A(cpuregs_13_[25]), .B(decoded_rs1_1_bF_buf31_), .C(decoded_rs1_0_bF_buf55_), .Y(_9555_) );
AOI21X1 AOI21X1_622 ( .A(_7128_), .B(decoded_rs1_1_bF_buf30_), .C(_9555_), .Y(_9556_) );
NOR2X1 NOR2X1_824 ( .A(cpuregs_14_[25]), .B(_7556__bF_buf31), .Y(_9557_) );
OAI21X1 OAI21X1_1965 ( .A(cpuregs_12_[25]), .B(decoded_rs1_1_bF_buf29_), .C(_7569__bF_buf21), .Y(_9558_) );
OAI21X1 OAI21X1_1966 ( .A(_9557_), .B(_9558_), .C(decoded_rs1_2_bF_buf10_), .Y(_9559_) );
OAI22X1 OAI22X1_192 ( .A(_9554_), .B(_9551_), .C(_9556_), .D(_9559_), .Y(_9560_) );
NAND2X1 NAND2X1_586 ( .A(_7552__bF_buf4), .B(_9560_), .Y(_9561_) );
OAI21X1 OAI21X1_1967 ( .A(_9548_), .B(_7552__bF_buf3), .C(_9561_), .Y(_9562_) );
NAND2X1 NAND2X1_587 ( .A(decoded_rs1_3_bF_buf1_), .B(_9562_), .Y(_9563_) );
AND2X2 AND2X2_127 ( .A(cpuregs_17_[25]), .B(decoded_rs1_0_bF_buf54_), .Y(_9564_) );
OAI21X1 OAI21X1_1968 ( .A(_7150_), .B(decoded_rs1_0_bF_buf53_), .C(_7556__bF_buf30), .Y(_9565_) );
AND2X2 AND2X2_128 ( .A(_7569__bF_buf20), .B(cpuregs_18_[25]), .Y(_9566_) );
OAI21X1 OAI21X1_1969 ( .A(_7153_), .B(_7569__bF_buf19), .C(decoded_rs1_1_bF_buf28_), .Y(_9567_) );
OAI22X1 OAI22X1_193 ( .A(_9565_), .B(_9564_), .C(_9567_), .D(_9566_), .Y(_9568_) );
INVX1 INVX1_800 ( .A(cpuregs_21_[25]), .Y(_9569_) );
AOI21X1 AOI21X1_623 ( .A(cpuregs_20_[25]), .B(_7569__bF_buf18), .C(decoded_rs1_1_bF_buf27_), .Y(_9570_) );
OAI21X1 OAI21X1_1970 ( .A(_9569_), .B(_7569__bF_buf17), .C(_9570_), .Y(_9571_) );
AOI21X1 AOI21X1_624 ( .A(cpuregs_23_[25]), .B(decoded_rs1_0_bF_buf52_), .C(_7556__bF_buf29), .Y(_9572_) );
OAI21X1 OAI21X1_1971 ( .A(_7161_), .B(decoded_rs1_0_bF_buf51_), .C(_9572_), .Y(_9573_) );
NAND3X1 NAND3X1_48 ( .A(decoded_rs1_2_bF_buf9_), .B(_9571_), .C(_9573_), .Y(_9574_) );
OAI21X1 OAI21X1_1972 ( .A(decoded_rs1_2_bF_buf8_), .B(_9568_), .C(_9574_), .Y(_9575_) );
NOR2X1 NOR2X1_825 ( .A(cpuregs_1_[25]), .B(decoded_rs1_2_bF_buf7_), .Y(_9576_) );
OAI21X1 OAI21X1_1973 ( .A(_7560__bF_buf11), .B(cpuregs_5_[25]), .C(decoded_rs1_0_bF_buf50_), .Y(_9577_) );
OAI21X1 OAI21X1_1974 ( .A(_7560__bF_buf10), .B(cpuregs_4_[25]), .C(_7569__bF_buf16), .Y(_9578_) );
AOI21X1 AOI21X1_625 ( .A(_7105_), .B(_7560__bF_buf9), .C(_9578_), .Y(_9579_) );
NOR2X1 NOR2X1_826 ( .A(decoded_rs1_1_bF_buf26_), .B(_9579_), .Y(_9580_) );
OAI21X1 OAI21X1_1975 ( .A(_9576_), .B(_9577_), .C(_9580_), .Y(_9581_) );
NOR2X1 NOR2X1_827 ( .A(cpuregs_3_[25]), .B(decoded_rs1_2_bF_buf6_), .Y(_9582_) );
OAI21X1 OAI21X1_1976 ( .A(_7560__bF_buf8), .B(cpuregs_7_[25]), .C(decoded_rs1_0_bF_buf49_), .Y(_9583_) );
NOR2X1 NOR2X1_828 ( .A(_9582_), .B(_9583_), .Y(_9584_) );
NOR2X1 NOR2X1_829 ( .A(cpuregs_2_[25]), .B(decoded_rs1_2_bF_buf5_), .Y(_9585_) );
OAI21X1 OAI21X1_1977 ( .A(_7560__bF_buf7), .B(cpuregs_6_[25]), .C(_7569__bF_buf15), .Y(_9586_) );
OAI21X1 OAI21X1_1978 ( .A(_9586_), .B(_9585_), .C(decoded_rs1_1_bF_buf25_), .Y(_9587_) );
OAI21X1 OAI21X1_1979 ( .A(_9584_), .B(_9587_), .C(_9581_), .Y(_9588_) );
NAND2X1 NAND2X1_588 ( .A(_7552__bF_buf2), .B(_9588_), .Y(_9589_) );
OAI21X1 OAI21X1_1980 ( .A(_7552__bF_buf1), .B(_9575_), .C(_9589_), .Y(_9590_) );
AOI21X1 AOI21X1_626 ( .A(_7561__bF_buf4), .B(_9590_), .C(_7586__bF_buf2), .Y(_9591_) );
AOI22X1 AOI22X1_94 ( .A(reg_pc_25_), .B(_7551__bF_buf3), .C(_9591_), .D(_9563_), .Y(_9592_) );
OAI21X1 OAI21X1_1981 ( .A(instr_slli), .B(instr_sll), .C(_10734__24_), .Y(_9593_) );
OAI21X1 OAI21X1_1982 ( .A(_7698__bF_buf1), .B(_5021_), .C(_9593_), .Y(_9594_) );
AND2X2 AND2X2_129 ( .A(_9594_), .B(_4579__bF_buf3), .Y(_9595_) );
OAI21X1 OAI21X1_1983 ( .A(_7778_), .B(_7700__bF_buf4), .C(_10734__29_), .Y(_9596_) );
AOI21X1 AOI21X1_627 ( .A(_9343_), .B(_9596_), .C(_4579__bF_buf2), .Y(_9597_) );
OAI21X1 OAI21X1_1984 ( .A(_9595_), .B(_9597_), .C(_4584_), .Y(_9598_) );
OAI21X1 OAI21X1_1985 ( .A(_7627_), .B(_5027_), .C(resetn_bF_buf10), .Y(_9599_) );
AOI21X1 AOI21X1_628 ( .A(_10734__25_), .B(_4597__bF_buf1), .C(_9599_), .Y(_9600_) );
AND2X2 AND2X2_130 ( .A(_9598_), .B(_9600_), .Y(_9601_) );
OAI21X1 OAI21X1_1986 ( .A(_9592_), .B(_4538__bF_buf0), .C(_9601_), .Y(_9602_) );
AOI21X1 AOI21X1_629 ( .A(_9537_), .B(_9536_), .C(_9602_), .Y(_9603_) );
AOI22X1 AOI22X1_95 ( .A(_4426__bF_buf5), .B(_5027_), .C(_9603_), .D(_9535_), .Y(_81__25_) );
NOR2X1 NOR2X1_830 ( .A(_9521_), .B(_9526_), .Y(_9604_) );
INVX1 INVX1_801 ( .A(_9604_), .Y(_9605_) );
NOR2X1 NOR2X1_831 ( .A(_10734__26_), .B(decoded_imm_26_), .Y(_9606_) );
INVX1 INVX1_802 ( .A(decoded_imm_26_), .Y(_9607_) );
NOR2X1 NOR2X1_832 ( .A(_5021_), .B(_9607_), .Y(_9608_) );
NOR2X1 NOR2X1_833 ( .A(_9606_), .B(_9608_), .Y(_9609_) );
OAI21X1 OAI21X1_1987 ( .A(_9531_), .B(_9605_), .C(_9609_), .Y(_9610_) );
NOR2X1 NOR2X1_834 ( .A(_9605_), .B(_9531_), .Y(_9611_) );
OAI21X1 OAI21X1_1988 ( .A(_9606_), .B(_9608_), .C(_9611_), .Y(_9612_) );
AND2X2 AND2X2_131 ( .A(_9612_), .B(_9610_), .Y(_9613_) );
AOI21X1 AOI21X1_630 ( .A(_5021_), .B(_7631__bF_buf1), .C(_7629__bF_buf2), .Y(_9614_) );
OAI21X1 OAI21X1_1989 ( .A(_9613_), .B(_7631__bF_buf0), .C(_9614_), .Y(_9615_) );
AOI21X1 AOI21X1_631 ( .A(_5021_), .B(_7623__bF_buf0), .C(_4587__bF_buf1), .Y(_9616_) );
OAI21X1 OAI21X1_1990 ( .A(_9613_), .B(_7623__bF_buf4), .C(_9616_), .Y(_9617_) );
OAI21X1 OAI21X1_1991 ( .A(_7201_), .B(decoded_rs1_0_bF_buf48_), .C(_7556__bF_buf28), .Y(_9618_) );
AOI21X1 AOI21X1_632 ( .A(cpuregs_25_[26]), .B(decoded_rs1_0_bF_buf47_), .C(_9618_), .Y(_9619_) );
NAND2X1 NAND2X1_589 ( .A(_7197_), .B(_7569__bF_buf14), .Y(_9620_) );
OAI21X1 OAI21X1_1992 ( .A(cpuregs_27_[26]), .B(_7569__bF_buf13), .C(_9620_), .Y(_9621_) );
AOI21X1 AOI21X1_633 ( .A(decoded_rs1_1_bF_buf24_), .B(_9621_), .C(_9619_), .Y(_9622_) );
NOR2X1 NOR2X1_835 ( .A(_7209_), .B(_7569__bF_buf12), .Y(_9623_) );
OAI21X1 OAI21X1_1993 ( .A(_7207_), .B(decoded_rs1_0_bF_buf46_), .C(_7556__bF_buf27), .Y(_9624_) );
AOI21X1 AOI21X1_634 ( .A(cpuregs_31_[26]), .B(decoded_rs1_0_bF_buf45_), .C(_7556__bF_buf26), .Y(_9625_) );
OAI21X1 OAI21X1_1994 ( .A(_7204_), .B(decoded_rs1_0_bF_buf44_), .C(_9625_), .Y(_9626_) );
OAI21X1 OAI21X1_1995 ( .A(_9623_), .B(_9624_), .C(_9626_), .Y(_9627_) );
OAI21X1 OAI21X1_1996 ( .A(_9627_), .B(_7560__bF_buf6), .C(decoded_rs1_3_bF_buf0_), .Y(_9628_) );
AOI21X1 AOI21X1_635 ( .A(_7560__bF_buf5), .B(_9622_), .C(_9628_), .Y(_9629_) );
MUX2X1 MUX2X1_190 ( .A(cpuregs_18_[26]), .B(cpuregs_16_[26]), .S(decoded_rs1_1_bF_buf23_), .Y(_9630_) );
NOR2X1 NOR2X1_836 ( .A(decoded_rs1_0_bF_buf43_), .B(_9630_), .Y(_9631_) );
MUX2X1 MUX2X1_191 ( .A(cpuregs_19_[26]), .B(cpuregs_17_[26]), .S(decoded_rs1_1_bF_buf22_), .Y(_9632_) );
OAI21X1 OAI21X1_1997 ( .A(_9632_), .B(_7569__bF_buf11), .C(_7560__bF_buf4), .Y(_9633_) );
OAI21X1 OAI21X1_1998 ( .A(_7221_), .B(decoded_rs1_0_bF_buf42_), .C(_7556__bF_buf25), .Y(_9634_) );
AOI21X1 AOI21X1_636 ( .A(cpuregs_21_[26]), .B(decoded_rs1_0_bF_buf41_), .C(_9634_), .Y(_9635_) );
NAND2X1 NAND2X1_590 ( .A(_7224_), .B(_7569__bF_buf10), .Y(_9636_) );
OAI21X1 OAI21X1_1999 ( .A(cpuregs_23_[26]), .B(_7569__bF_buf9), .C(_9636_), .Y(_9637_) );
AOI21X1 AOI21X1_637 ( .A(decoded_rs1_1_bF_buf21_), .B(_9637_), .C(_9635_), .Y(_9638_) );
OAI22X1 OAI22X1_194 ( .A(_9631_), .B(_9633_), .C(_9638_), .D(_7560__bF_buf3), .Y(_9639_) );
AND2X2 AND2X2_132 ( .A(_9639_), .B(_7561__bF_buf3), .Y(_9640_) );
OAI21X1 OAI21X1_2000 ( .A(_9640_), .B(_9629_), .C(decoded_rs1_4_bF_buf2_), .Y(_9641_) );
NOR2X1 NOR2X1_837 ( .A(_7183_), .B(_7569__bF_buf8), .Y(_9642_) );
INVX1 INVX1_803 ( .A(cpuregs_12_[26]), .Y(_9643_) );
OAI21X1 OAI21X1_2001 ( .A(_9643_), .B(decoded_rs1_0_bF_buf40_), .C(_7556__bF_buf24), .Y(_9644_) );
AND2X2 AND2X2_133 ( .A(_7569__bF_buf7), .B(cpuregs_14_[26]), .Y(_9645_) );
INVX1 INVX1_804 ( .A(cpuregs_15_[26]), .Y(_9646_) );
OAI21X1 OAI21X1_2002 ( .A(_9646_), .B(_7569__bF_buf6), .C(decoded_rs1_1_bF_buf20_), .Y(_9647_) );
OAI22X1 OAI22X1_195 ( .A(_9644_), .B(_9642_), .C(_9647_), .D(_9645_), .Y(_9648_) );
MUX2X1 MUX2X1_192 ( .A(cpuregs_9_[26]), .B(cpuregs_8_[26]), .S(decoded_rs1_0_bF_buf39_), .Y(_9649_) );
MUX2X1 MUX2X1_193 ( .A(cpuregs_11_[26]), .B(cpuregs_10_[26]), .S(decoded_rs1_0_bF_buf38_), .Y(_9650_) );
MUX2X1 MUX2X1_194 ( .A(_9650_), .B(_9649_), .S(decoded_rs1_1_bF_buf19_), .Y(_9651_) );
AOI21X1 AOI21X1_638 ( .A(_7560__bF_buf2), .B(_9651_), .C(_7561__bF_buf2), .Y(_9652_) );
OAI21X1 OAI21X1_2003 ( .A(_7560__bF_buf1), .B(_9648_), .C(_9652_), .Y(_9653_) );
OAI21X1 OAI21X1_2004 ( .A(_7560__bF_buf0), .B(cpuregs_5_[26]), .C(decoded_rs1_0_bF_buf37_), .Y(_9654_) );
AOI21X1 AOI21X1_639 ( .A(_7170_), .B(_7560__bF_buf12), .C(_9654_), .Y(_9655_) );
NOR2X1 NOR2X1_838 ( .A(cpuregs_0_[26]), .B(decoded_rs1_2_bF_buf4_), .Y(_9656_) );
OAI21X1 OAI21X1_2005 ( .A(_7560__bF_buf11), .B(cpuregs_4_[26]), .C(_7569__bF_buf5), .Y(_9657_) );
OAI21X1 OAI21X1_2006 ( .A(_9657_), .B(_9656_), .C(_7556__bF_buf23), .Y(_9658_) );
NOR2X1 NOR2X1_839 ( .A(_9655_), .B(_9658_), .Y(_9659_) );
NOR2X1 NOR2X1_840 ( .A(cpuregs_3_[26]), .B(decoded_rs1_2_bF_buf3_), .Y(_9660_) );
OAI21X1 OAI21X1_2007 ( .A(_7560__bF_buf10), .B(cpuregs_7_[26]), .C(decoded_rs1_0_bF_buf36_), .Y(_9661_) );
NOR2X1 NOR2X1_841 ( .A(_9660_), .B(_9661_), .Y(_9662_) );
NOR2X1 NOR2X1_842 ( .A(cpuregs_2_[26]), .B(decoded_rs1_2_bF_buf2_), .Y(_9663_) );
OAI21X1 OAI21X1_2008 ( .A(_7560__bF_buf9), .B(cpuregs_6_[26]), .C(_7569__bF_buf4), .Y(_9664_) );
OAI21X1 OAI21X1_2009 ( .A(_9664_), .B(_9663_), .C(decoded_rs1_1_bF_buf18_), .Y(_9665_) );
NOR2X1 NOR2X1_843 ( .A(_9662_), .B(_9665_), .Y(_9666_) );
OAI21X1 OAI21X1_2010 ( .A(_9659_), .B(_9666_), .C(_7561__bF_buf1), .Y(_9667_) );
NAND2X1 NAND2X1_591 ( .A(_9653_), .B(_9667_), .Y(_9668_) );
AOI21X1 AOI21X1_640 ( .A(_7552__bF_buf0), .B(_9668_), .C(_7586__bF_buf1), .Y(_9669_) );
NAND2X1 NAND2X1_592 ( .A(_9669_), .B(_9641_), .Y(_9670_) );
OAI21X1 OAI21X1_2011 ( .A(_4860_), .B(_7643_), .C(_9670_), .Y(_9671_) );
INVX1 INVX1_805 ( .A(_9420_), .Y(_9672_) );
OAI21X1 OAI21X1_2012 ( .A(_7698__bF_buf0), .B(_4998_), .C(_4580__bF_buf3), .Y(_9673_) );
OAI21X1 OAI21X1_2013 ( .A(_5027_), .B(_7700__bF_buf3), .C(_4579__bF_buf1), .Y(_9674_) );
OAI22X1 OAI22X1_196 ( .A(_9423_), .B(_9674_), .C(_9673_), .D(_9672_), .Y(_9675_) );
OAI21X1 OAI21X1_2014 ( .A(_7627_), .B(_5021_), .C(resetn_bF_buf9), .Y(_9676_) );
AOI21X1 AOI21X1_641 ( .A(_10734__26_), .B(_4597__bF_buf0), .C(_9676_), .Y(_9677_) );
OAI21X1 OAI21X1_2015 ( .A(_7697__bF_buf3), .B(_9675_), .C(_9677_), .Y(_9678_) );
AOI21X1 AOI21X1_642 ( .A(cpu_state_2_bF_buf4_), .B(_9671_), .C(_9678_), .Y(_9679_) );
AND2X2 AND2X2_134 ( .A(_9617_), .B(_9679_), .Y(_9680_) );
AOI22X1 AOI22X1_96 ( .A(_4426__bF_buf4), .B(_5021_), .C(_9680_), .D(_9615_), .Y(_81__26_) );
OAI21X1 OAI21X1_2016 ( .A(_5021_), .B(_9607_), .C(_9610_), .Y(_9681_) );
NOR2X1 NOR2X1_844 ( .A(_10734__27_), .B(decoded_imm_27_), .Y(_9682_) );
INVX1 INVX1_806 ( .A(decoded_imm_27_), .Y(_9683_) );
NOR2X1 NOR2X1_845 ( .A(_5016_), .B(_9683_), .Y(_9684_) );
NOR2X1 NOR2X1_846 ( .A(_9682_), .B(_9684_), .Y(_9685_) );
INVX1 INVX1_807 ( .A(_9685_), .Y(_9686_) );
OR2X2 OR2X2_16 ( .A(_9681_), .B(_9686_), .Y(_9687_) );
OAI21X1 OAI21X1_2017 ( .A(_9682_), .B(_9684_), .C(_9681_), .Y(_9688_) );
NAND2X1 NAND2X1_593 ( .A(_9688_), .B(_9687_), .Y(_9689_) );
AOI21X1 AOI21X1_643 ( .A(_5016_), .B(_7631__bF_buf5), .C(_7629__bF_buf1), .Y(_9690_) );
OAI21X1 OAI21X1_2018 ( .A(_9689_), .B(_7631__bF_buf4), .C(_9690_), .Y(_9691_) );
NAND3X1 NAND3X1_49 ( .A(_7624__bF_buf2), .B(_9688_), .C(_9687_), .Y(_9692_) );
AOI21X1 AOI21X1_644 ( .A(_5016_), .B(_7623__bF_buf3), .C(_4587__bF_buf0), .Y(_9693_) );
AND2X2 AND2X2_135 ( .A(cpuregs_17_[27]), .B(decoded_rs1_0_bF_buf35_), .Y(_9694_) );
OAI21X1 OAI21X1_2019 ( .A(_7277_), .B(decoded_rs1_0_bF_buf34_), .C(_7556__bF_buf22), .Y(_9695_) );
AND2X2 AND2X2_136 ( .A(_7569__bF_buf3), .B(cpuregs_18_[27]), .Y(_9696_) );
OAI21X1 OAI21X1_2020 ( .A(_7280_), .B(_7569__bF_buf2), .C(decoded_rs1_1_bF_buf17_), .Y(_9697_) );
OAI22X1 OAI22X1_197 ( .A(_9695_), .B(_9694_), .C(_9697_), .D(_9696_), .Y(_9698_) );
NOR2X1 NOR2X1_847 ( .A(decoded_rs1_2_bF_buf1_), .B(_9698_), .Y(_9699_) );
AND2X2 AND2X2_137 ( .A(cpuregs_21_[27]), .B(decoded_rs1_0_bF_buf33_), .Y(_9700_) );
OAI21X1 OAI21X1_2021 ( .A(_7285_), .B(decoded_rs1_0_bF_buf32_), .C(_7556__bF_buf21), .Y(_9701_) );
NOR2X1 NOR2X1_848 ( .A(decoded_rs1_0_bF_buf31_), .B(_7288_), .Y(_9702_) );
INVX1 INVX1_808 ( .A(cpuregs_23_[27]), .Y(_9703_) );
OAI21X1 OAI21X1_2022 ( .A(_9703_), .B(_7569__bF_buf1), .C(decoded_rs1_1_bF_buf16_), .Y(_9704_) );
OAI22X1 OAI22X1_198 ( .A(_9701_), .B(_9700_), .C(_9704_), .D(_9702_), .Y(_9705_) );
OAI21X1 OAI21X1_2023 ( .A(_9705_), .B(_7560__bF_buf8), .C(_7561__bF_buf0), .Y(_9706_) );
NOR2X1 NOR2X1_849 ( .A(_9699_), .B(_9706_), .Y(_9707_) );
AOI21X1 AOI21X1_645 ( .A(_7269_), .B(_7556__bF_buf20), .C(decoded_rs1_0_bF_buf30_), .Y(_9708_) );
OAI21X1 OAI21X1_2024 ( .A(cpuregs_30_[27]), .B(_7556__bF_buf19), .C(_9708_), .Y(_9709_) );
NOR2X1 NOR2X1_850 ( .A(cpuregs_31_[27]), .B(_7556__bF_buf18), .Y(_9710_) );
OAI21X1 OAI21X1_2025 ( .A(cpuregs_29_[27]), .B(decoded_rs1_1_bF_buf15_), .C(decoded_rs1_0_bF_buf29_), .Y(_9711_) );
OAI21X1 OAI21X1_2026 ( .A(_9710_), .B(_9711_), .C(_9709_), .Y(_9712_) );
OAI21X1 OAI21X1_2027 ( .A(cpuregs_24_[27]), .B(decoded_rs1_1_bF_buf14_), .C(_7569__bF_buf0), .Y(_9713_) );
AOI21X1 AOI21X1_646 ( .A(_7262_), .B(decoded_rs1_1_bF_buf13_), .C(_9713_), .Y(_9714_) );
INVX1 INVX1_809 ( .A(cpuregs_27_[27]), .Y(_9715_) );
OAI21X1 OAI21X1_2028 ( .A(cpuregs_25_[27]), .B(decoded_rs1_1_bF_buf12_), .C(decoded_rs1_0_bF_buf28_), .Y(_9716_) );
AOI21X1 AOI21X1_647 ( .A(_9715_), .B(decoded_rs1_1_bF_buf11_), .C(_9716_), .Y(_9717_) );
OAI21X1 OAI21X1_2029 ( .A(_9714_), .B(_9717_), .C(_7560__bF_buf7), .Y(_9718_) );
NAND2X1 NAND2X1_594 ( .A(decoded_rs1_3_bF_buf6_), .B(_9718_), .Y(_9719_) );
AOI21X1 AOI21X1_648 ( .A(decoded_rs1_2_bF_buf0_), .B(_9712_), .C(_9719_), .Y(_9720_) );
OAI21X1 OAI21X1_2030 ( .A(_9720_), .B(_9707_), .C(decoded_rs1_4_bF_buf1_), .Y(_9721_) );
INVX1 INVX1_810 ( .A(cpuregs_12_[27]), .Y(_9722_) );
AOI21X1 AOI21X1_649 ( .A(_9722_), .B(_7556__bF_buf17), .C(decoded_rs1_0_bF_buf27_), .Y(_9723_) );
OAI21X1 OAI21X1_2031 ( .A(cpuregs_14_[27]), .B(_7556__bF_buf16), .C(_9723_), .Y(_9724_) );
AOI21X1 AOI21X1_650 ( .A(_7247_), .B(_7556__bF_buf15), .C(_7569__bF_buf48), .Y(_9725_) );
OAI21X1 OAI21X1_2032 ( .A(cpuregs_15_[27]), .B(_7556__bF_buf14), .C(_9725_), .Y(_9726_) );
AOI21X1 AOI21X1_651 ( .A(_9724_), .B(_9726_), .C(_7560__bF_buf6), .Y(_9727_) );
AND2X2 AND2X2_138 ( .A(cpuregs_1_[27]), .B(decoded_rs1_0_bF_buf26_), .Y(_9728_) );
INVX1 INVX1_811 ( .A(cpuregs_0_[27]), .Y(_9729_) );
OAI21X1 OAI21X1_2033 ( .A(_9729_), .B(decoded_rs1_0_bF_buf25_), .C(_7556__bF_buf13), .Y(_9730_) );
NOR2X1 NOR2X1_851 ( .A(decoded_rs1_0_bF_buf24_), .B(_7233_), .Y(_9731_) );
INVX1 INVX1_812 ( .A(cpuregs_3_[27]), .Y(_9732_) );
OAI21X1 OAI21X1_2034 ( .A(_9732_), .B(_7569__bF_buf47), .C(decoded_rs1_1_bF_buf10_), .Y(_9733_) );
OAI22X1 OAI22X1_199 ( .A(_9730_), .B(_9728_), .C(_9733_), .D(_9731_), .Y(_9734_) );
NOR2X1 NOR2X1_852 ( .A(decoded_rs1_2_bF_buf12_), .B(_9734_), .Y(_9735_) );
AND2X2 AND2X2_139 ( .A(cpuregs_5_[27]), .B(decoded_rs1_0_bF_buf23_), .Y(_9736_) );
INVX1 INVX1_813 ( .A(cpuregs_4_[27]), .Y(_9737_) );
OAI21X1 OAI21X1_2035 ( .A(_9737_), .B(decoded_rs1_0_bF_buf22_), .C(_7556__bF_buf12), .Y(_9738_) );
NOR2X1 NOR2X1_853 ( .A(decoded_rs1_0_bF_buf21_), .B(_7240_), .Y(_9739_) );
INVX1 INVX1_814 ( .A(cpuregs_7_[27]), .Y(_9740_) );
OAI21X1 OAI21X1_2036 ( .A(_9740_), .B(_7569__bF_buf46), .C(decoded_rs1_1_bF_buf9_), .Y(_9741_) );
OAI22X1 OAI22X1_200 ( .A(_9738_), .B(_9736_), .C(_9741_), .D(_9739_), .Y(_9742_) );
OAI21X1 OAI21X1_2037 ( .A(_9742_), .B(_7560__bF_buf5), .C(_7561__bF_buf6), .Y(_9743_) );
INVX1 INVX1_815 ( .A(cpuregs_8_[27]), .Y(_9744_) );
AOI21X1 AOI21X1_652 ( .A(_9744_), .B(_7556__bF_buf11), .C(decoded_rs1_0_bF_buf20_), .Y(_9745_) );
OAI21X1 OAI21X1_2038 ( .A(cpuregs_10_[27]), .B(_7556__bF_buf10), .C(_9745_), .Y(_9746_) );
AOI21X1 AOI21X1_653 ( .A(_7254_), .B(_7556__bF_buf9), .C(_7569__bF_buf45), .Y(_9747_) );
OAI21X1 OAI21X1_2039 ( .A(cpuregs_11_[27]), .B(_7556__bF_buf8), .C(_9747_), .Y(_9748_) );
AND2X2 AND2X2_140 ( .A(_9746_), .B(_9748_), .Y(_9749_) );
OAI21X1 OAI21X1_2040 ( .A(_9749_), .B(decoded_rs1_2_bF_buf11_), .C(decoded_rs1_3_bF_buf5_), .Y(_9750_) );
OAI22X1 OAI22X1_201 ( .A(_9735_), .B(_9743_), .C(_9750_), .D(_9727_), .Y(_9751_) );
AOI21X1 AOI21X1_654 ( .A(_7552__bF_buf5), .B(_9751_), .C(_7586__bF_buf0), .Y(_9752_) );
AOI22X1 AOI22X1_97 ( .A(reg_pc_27_), .B(_7551__bF_buf2), .C(_9752_), .D(_9721_), .Y(_9753_) );
NOR2X1 NOR2X1_854 ( .A(_4538__bF_buf4), .B(_9753_), .Y(_9754_) );
OAI21X1 OAI21X1_2041 ( .A(instr_slli), .B(instr_sll), .C(_10734__26_), .Y(_9755_) );
OAI21X1 OAI21X1_2042 ( .A(_7698__bF_buf4), .B(_5004_), .C(_9755_), .Y(_9756_) );
OAI21X1 OAI21X1_2043 ( .A(_7698__bF_buf3), .B(_4991_), .C(_9510_), .Y(_9757_) );
MUX2X1 MUX2X1_195 ( .A(_9756_), .B(_9757_), .S(_4579__bF_buf0), .Y(_9758_) );
OAI21X1 OAI21X1_2044 ( .A(_7627_), .B(_5016_), .C(resetn_bF_buf8), .Y(_9759_) );
AOI21X1 AOI21X1_655 ( .A(_10734__27_), .B(_4597__bF_buf3), .C(_9759_), .Y(_9760_) );
OAI21X1 OAI21X1_2045 ( .A(_7697__bF_buf2), .B(_9758_), .C(_9760_), .Y(_9761_) );
OR2X2 OR2X2_17 ( .A(_9754_), .B(_9761_), .Y(_9762_) );
AOI21X1 AOI21X1_656 ( .A(_9693_), .B(_9692_), .C(_9762_), .Y(_9763_) );
AOI22X1 AOI22X1_98 ( .A(_4426__bF_buf3), .B(_5016_), .C(_9763_), .D(_9691_), .Y(_81__27_) );
NAND2X1 NAND2X1_595 ( .A(_9685_), .B(_9609_), .Y(_9764_) );
OR2X2 OR2X2_18 ( .A(_9530_), .B(_9764_), .Y(_9765_) );
AOI21X1 AOI21X1_657 ( .A(_9436_), .B(_9528_), .C(_9765_), .Y(_9766_) );
AOI21X1 AOI21X1_658 ( .A(_9608_), .B(_9685_), .C(_9684_), .Y(_9767_) );
OAI21X1 OAI21X1_2046 ( .A(_9604_), .B(_9764_), .C(_9767_), .Y(_9768_) );
NOR2X1 NOR2X1_855 ( .A(_10734__28_), .B(decoded_imm_28_), .Y(_9769_) );
INVX1 INVX1_816 ( .A(decoded_imm_28_), .Y(_9770_) );
NOR2X1 NOR2X1_856 ( .A(_5004_), .B(_9770_), .Y(_9771_) );
NOR2X1 NOR2X1_857 ( .A(_9769_), .B(_9771_), .Y(_9772_) );
OAI21X1 OAI21X1_2047 ( .A(_9766_), .B(_9768_), .C(_9772_), .Y(_9773_) );
INVX1 INVX1_817 ( .A(_9765_), .Y(_9774_) );
AOI21X1 AOI21X1_659 ( .A(_9774_), .B(_9439_), .C(_9768_), .Y(_9775_) );
OAI21X1 OAI21X1_2048 ( .A(_9769_), .B(_9771_), .C(_9775_), .Y(_9776_) );
NAND2X1 NAND2X1_596 ( .A(_9773_), .B(_9776_), .Y(_9777_) );
OAI21X1 OAI21X1_2049 ( .A(_7632__bF_buf1), .B(_10734__28_), .C(_7630_), .Y(_9778_) );
AOI21X1 AOI21X1_660 ( .A(_7632__bF_buf0), .B(_9777_), .C(_9778_), .Y(_9779_) );
NAND2X1 NAND2X1_597 ( .A(_7624__bF_buf1), .B(_9777_), .Y(_9780_) );
AOI21X1 AOI21X1_661 ( .A(_5004_), .B(_7623__bF_buf2), .C(_4587__bF_buf3), .Y(_9781_) );
NAND2X1 NAND2X1_598 ( .A(_9781_), .B(_9780_), .Y(_9782_) );
AND2X2 AND2X2_141 ( .A(cpuregs_17_[28]), .B(decoded_rs1_0_bF_buf19_), .Y(_9783_) );
INVX1 INVX1_818 ( .A(cpuregs_16_[28]), .Y(_9784_) );
OAI21X1 OAI21X1_2050 ( .A(_9784_), .B(decoded_rs1_0_bF_buf18_), .C(_7556__bF_buf7), .Y(_9785_) );
AND2X2 AND2X2_142 ( .A(_7569__bF_buf44), .B(cpuregs_18_[28]), .Y(_9786_) );
INVX1 INVX1_819 ( .A(cpuregs_19_[28]), .Y(_9787_) );
OAI21X1 OAI21X1_2051 ( .A(_9787_), .B(_7569__bF_buf43), .C(decoded_rs1_1_bF_buf8_), .Y(_9788_) );
OAI22X1 OAI22X1_202 ( .A(_9785_), .B(_9783_), .C(_9788_), .D(_9786_), .Y(_9789_) );
NOR2X1 NOR2X1_858 ( .A(decoded_rs1_2_bF_buf10_), .B(_9789_), .Y(_9790_) );
NOR2X1 NOR2X1_859 ( .A(_7300_), .B(_7569__bF_buf42), .Y(_9791_) );
OAI21X1 OAI21X1_2052 ( .A(_7297_), .B(decoded_rs1_0_bF_buf17_), .C(_7556__bF_buf6), .Y(_9792_) );
NOR2X1 NOR2X1_860 ( .A(decoded_rs1_0_bF_buf16_), .B(_7304_), .Y(_9793_) );
OAI21X1 OAI21X1_2053 ( .A(_7307_), .B(_7569__bF_buf41), .C(decoded_rs1_1_bF_buf7_), .Y(_9794_) );
OAI22X1 OAI22X1_203 ( .A(_9792_), .B(_9791_), .C(_9794_), .D(_9793_), .Y(_9795_) );
OAI21X1 OAI21X1_2054 ( .A(_9795_), .B(_7560__bF_buf4), .C(_7561__bF_buf5), .Y(_9796_) );
NOR2X1 NOR2X1_861 ( .A(_9790_), .B(_9796_), .Y(_9797_) );
AOI21X1 AOI21X1_662 ( .A(_7335_), .B(_7556__bF_buf5), .C(decoded_rs1_0_bF_buf15_), .Y(_9798_) );
OAI21X1 OAI21X1_2055 ( .A(cpuregs_26_[28]), .B(_7556__bF_buf4), .C(_9798_), .Y(_9799_) );
NOR2X1 NOR2X1_862 ( .A(cpuregs_27_[28]), .B(_7556__bF_buf3), .Y(_9800_) );
OAI21X1 OAI21X1_2056 ( .A(cpuregs_25_[28]), .B(decoded_rs1_1_bF_buf6_), .C(decoded_rs1_0_bF_buf14_), .Y(_9801_) );
OAI21X1 OAI21X1_2057 ( .A(_9800_), .B(_9801_), .C(_9799_), .Y(_9802_) );
INVX1 INVX1_820 ( .A(cpuregs_30_[28]), .Y(_9803_) );
OAI21X1 OAI21X1_2058 ( .A(cpuregs_28_[28]), .B(decoded_rs1_1_bF_buf5_), .C(_7569__bF_buf40), .Y(_9804_) );
AOI21X1 AOI21X1_663 ( .A(_9803_), .B(decoded_rs1_1_bF_buf4_), .C(_9804_), .Y(_9805_) );
OAI21X1 OAI21X1_2059 ( .A(cpuregs_29_[28]), .B(decoded_rs1_1_bF_buf3_), .C(decoded_rs1_0_bF_buf13_), .Y(_9806_) );
AOI21X1 AOI21X1_664 ( .A(_7330_), .B(decoded_rs1_1_bF_buf2_), .C(_9806_), .Y(_9807_) );
OAI21X1 OAI21X1_2060 ( .A(_9805_), .B(_9807_), .C(decoded_rs1_2_bF_buf9_), .Y(_9808_) );
NAND2X1 NAND2X1_599 ( .A(decoded_rs1_3_bF_buf4_), .B(_9808_), .Y(_9809_) );
AOI21X1 AOI21X1_665 ( .A(_7560__bF_buf3), .B(_9802_), .C(_9809_), .Y(_9810_) );
OAI21X1 OAI21X1_2061 ( .A(_9810_), .B(_9797_), .C(decoded_rs1_4_bF_buf0_), .Y(_9811_) );
INVX1 INVX1_821 ( .A(cpuregs_14_[28]), .Y(_9812_) );
OAI21X1 OAI21X1_2062 ( .A(cpuregs_12_[28]), .B(decoded_rs1_1_bF_buf1_), .C(_7569__bF_buf39), .Y(_9813_) );
AOI21X1 AOI21X1_666 ( .A(_9812_), .B(decoded_rs1_1_bF_buf0_), .C(_9813_), .Y(_9814_) );
INVX1 INVX1_822 ( .A(cpuregs_15_[28]), .Y(_9815_) );
OAI21X1 OAI21X1_2063 ( .A(cpuregs_13_[28]), .B(decoded_rs1_1_bF_buf44_), .C(decoded_rs1_0_bF_buf12_), .Y(_9816_) );
AOI21X1 AOI21X1_667 ( .A(_9815_), .B(decoded_rs1_1_bF_buf43_), .C(_9816_), .Y(_9817_) );
OAI21X1 OAI21X1_2064 ( .A(_9814_), .B(_9817_), .C(decoded_rs1_2_bF_buf8_), .Y(_9818_) );
INVX1 INVX1_823 ( .A(cpuregs_10_[28]), .Y(_9819_) );
OAI21X1 OAI21X1_2065 ( .A(cpuregs_8_[28]), .B(decoded_rs1_1_bF_buf42_), .C(_7569__bF_buf38), .Y(_9820_) );
AOI21X1 AOI21X1_668 ( .A(_9819_), .B(decoded_rs1_1_bF_buf41_), .C(_9820_), .Y(_9821_) );
INVX1 INVX1_824 ( .A(cpuregs_11_[28]), .Y(_9822_) );
OAI21X1 OAI21X1_2066 ( .A(cpuregs_9_[28]), .B(decoded_rs1_1_bF_buf40_), .C(decoded_rs1_0_bF_buf11_), .Y(_9823_) );
AOI21X1 AOI21X1_669 ( .A(_9822_), .B(decoded_rs1_1_bF_buf39_), .C(_9823_), .Y(_9824_) );
OAI21X1 OAI21X1_2067 ( .A(_9821_), .B(_9824_), .C(_7560__bF_buf2), .Y(_9825_) );
NAND2X1 NAND2X1_600 ( .A(_9825_), .B(_9818_), .Y(_9826_) );
AND2X2 AND2X2_143 ( .A(cpuregs_1_[28]), .B(decoded_rs1_0_bF_buf10_), .Y(_9827_) );
INVX1 INVX1_825 ( .A(cpuregs_0_[28]), .Y(_9828_) );
OAI21X1 OAI21X1_2068 ( .A(_9828_), .B(decoded_rs1_0_bF_buf9_), .C(_7556__bF_buf2), .Y(_9829_) );
NOR2X1 NOR2X1_863 ( .A(decoded_rs1_0_bF_buf8_), .B(_7318_), .Y(_9830_) );
INVX1 INVX1_826 ( .A(cpuregs_3_[28]), .Y(_9831_) );
OAI21X1 OAI21X1_2069 ( .A(_9831_), .B(_7569__bF_buf37), .C(decoded_rs1_1_bF_buf38_), .Y(_9832_) );
OAI22X1 OAI22X1_204 ( .A(_9829_), .B(_9827_), .C(_9832_), .D(_9830_), .Y(_9833_) );
NOR2X1 NOR2X1_864 ( .A(decoded_rs1_2_bF_buf7_), .B(_9833_), .Y(_9834_) );
AND2X2 AND2X2_144 ( .A(cpuregs_5_[28]), .B(decoded_rs1_0_bF_buf7_), .Y(_9835_) );
INVX1 INVX1_827 ( .A(cpuregs_4_[28]), .Y(_9836_) );
OAI21X1 OAI21X1_2070 ( .A(_9836_), .B(decoded_rs1_0_bF_buf6_), .C(_7556__bF_buf1), .Y(_9837_) );
NOR2X1 NOR2X1_865 ( .A(decoded_rs1_0_bF_buf5_), .B(_7312_), .Y(_9838_) );
INVX1 INVX1_828 ( .A(cpuregs_7_[28]), .Y(_9839_) );
OAI21X1 OAI21X1_2071 ( .A(_9839_), .B(_7569__bF_buf36), .C(decoded_rs1_1_bF_buf37_), .Y(_9840_) );
OAI22X1 OAI22X1_205 ( .A(_9837_), .B(_9835_), .C(_9840_), .D(_9838_), .Y(_9841_) );
OAI21X1 OAI21X1_2072 ( .A(_9841_), .B(_7560__bF_buf1), .C(_7561__bF_buf4), .Y(_9842_) );
OAI22X1 OAI22X1_206 ( .A(_9834_), .B(_9842_), .C(_9826_), .D(_7561__bF_buf3), .Y(_9843_) );
AOI21X1 AOI21X1_670 ( .A(_7552__bF_buf4), .B(_9843_), .C(_7586__bF_buf3), .Y(_9844_) );
AOI22X1 AOI22X1_99 ( .A(reg_pc_28_), .B(_7551__bF_buf1), .C(_9844_), .D(_9811_), .Y(_9845_) );
OR2X2 OR2X2_19 ( .A(_9845_), .B(_4538__bF_buf3), .Y(_9846_) );
INVX1 INVX1_829 ( .A(_9593_), .Y(_9847_) );
NAND3X1 NAND3X1_50 ( .A(_10734__31_), .B(_7700__bF_buf2), .C(_7615_), .Y(_9848_) );
OAI21X1 OAI21X1_2073 ( .A(reg_sh_4_), .B(_4578_), .C(_9848_), .Y(_9849_) );
OAI21X1 OAI21X1_2074 ( .A(instr_slli), .B(instr_sll), .C(_10734__27_), .Y(_9850_) );
NAND3X1 NAND3X1_51 ( .A(_4579__bF_buf4), .B(_9850_), .C(_9596_), .Y(_9851_) );
OAI21X1 OAI21X1_2075 ( .A(_9849_), .B(_9847_), .C(_9851_), .Y(_9852_) );
MUX2X1 MUX2X1_196 ( .A(_9852_), .B(_5004_), .S(_4582_), .Y(_9853_) );
AOI22X1 AOI22X1_100 ( .A(_10734__28_), .B(_8855_), .C(_9853_), .D(cpu_state_4_), .Y(_9854_) );
NAND3X1 NAND3X1_52 ( .A(_9846_), .B(_9854_), .C(_9782_), .Y(_9855_) );
OAI21X1 OAI21X1_2076 ( .A(_9855_), .B(_9779_), .C(resetn_bF_buf7), .Y(_9856_) );
OAI21X1 OAI21X1_2077 ( .A(resetn_bF_buf6), .B(_5004_), .C(_9856_), .Y(_81__28_) );
OAI21X1 OAI21X1_2078 ( .A(_5004_), .B(_9770_), .C(_9773_), .Y(_9857_) );
NOR2X1 NOR2X1_866 ( .A(_10734__29_), .B(decoded_imm_29_), .Y(_9858_) );
INVX1 INVX1_830 ( .A(decoded_imm_29_), .Y(_9859_) );
NOR2X1 NOR2X1_867 ( .A(_5009_), .B(_9859_), .Y(_9860_) );
NOR2X1 NOR2X1_868 ( .A(_9858_), .B(_9860_), .Y(_9861_) );
INVX1 INVX1_831 ( .A(_9861_), .Y(_9862_) );
OR2X2 OR2X2_20 ( .A(_9857_), .B(_9862_), .Y(_9863_) );
OAI21X1 OAI21X1_2079 ( .A(_9858_), .B(_9860_), .C(_9857_), .Y(_9864_) );
NAND2X1 NAND2X1_601 ( .A(_9864_), .B(_9863_), .Y(_9865_) );
AOI21X1 AOI21X1_671 ( .A(_5009_), .B(_7631__bF_buf3), .C(_7629__bF_buf0), .Y(_9866_) );
OAI21X1 OAI21X1_2080 ( .A(_9865_), .B(_7631__bF_buf2), .C(_9866_), .Y(_9867_) );
NAND3X1 NAND3X1_53 ( .A(_7624__bF_buf0), .B(_9864_), .C(_9863_), .Y(_9868_) );
AOI21X1 AOI21X1_672 ( .A(_5009_), .B(_7623__bF_buf1), .C(_4587__bF_buf2), .Y(_9869_) );
AND2X2 AND2X2_145 ( .A(cpuregs_17_[29]), .B(decoded_rs1_0_bF_buf4_), .Y(_9870_) );
OAI21X1 OAI21X1_2081 ( .A(_7402_), .B(decoded_rs1_0_bF_buf3_), .C(_7556__bF_buf0), .Y(_9871_) );
AND2X2 AND2X2_146 ( .A(_7569__bF_buf35), .B(cpuregs_18_[29]), .Y(_9872_) );
OAI21X1 OAI21X1_2082 ( .A(_7405_), .B(_7569__bF_buf34), .C(decoded_rs1_1_bF_buf36_), .Y(_9873_) );
OAI22X1 OAI22X1_207 ( .A(_9871_), .B(_9870_), .C(_9873_), .D(_9872_), .Y(_9874_) );
NOR2X1 NOR2X1_869 ( .A(decoded_rs1_2_bF_buf6_), .B(_9874_), .Y(_9875_) );
AND2X2 AND2X2_147 ( .A(cpuregs_21_[29]), .B(decoded_rs1_0_bF_buf2_), .Y(_9876_) );
OAI21X1 OAI21X1_2083 ( .A(_7410_), .B(decoded_rs1_0_bF_buf1_), .C(_7556__bF_buf42), .Y(_9877_) );
NOR2X1 NOR2X1_870 ( .A(decoded_rs1_0_bF_buf0_), .B(_7413_), .Y(_9878_) );
INVX1 INVX1_832 ( .A(cpuregs_23_[29]), .Y(_9879_) );
OAI21X1 OAI21X1_2084 ( .A(_9879_), .B(_7569__bF_buf33), .C(decoded_rs1_1_bF_buf35_), .Y(_9880_) );
OAI22X1 OAI22X1_208 ( .A(_9877_), .B(_9876_), .C(_9880_), .D(_9878_), .Y(_9881_) );
OAI21X1 OAI21X1_2085 ( .A(_9881_), .B(_7560__bF_buf0), .C(_7561__bF_buf2), .Y(_9882_) );
NOR2X1 NOR2X1_871 ( .A(_9875_), .B(_9882_), .Y(_9883_) );
OAI21X1 OAI21X1_2086 ( .A(_7394_), .B(decoded_rs1_0_bF_buf57_), .C(_7556__bF_buf41), .Y(_9884_) );
AOI21X1 AOI21X1_673 ( .A(cpuregs_29_[29]), .B(decoded_rs1_0_bF_buf56_), .C(_9884_), .Y(_9885_) );
INVX1 INVX1_833 ( .A(cpuregs_31_[29]), .Y(_9886_) );
OAI21X1 OAI21X1_2087 ( .A(_9886_), .B(_7569__bF_buf32), .C(decoded_rs1_1_bF_buf34_), .Y(_9887_) );
AOI21X1 AOI21X1_674 ( .A(cpuregs_30_[29]), .B(_7569__bF_buf31), .C(_9887_), .Y(_9888_) );
OAI21X1 OAI21X1_2088 ( .A(_9888_), .B(_9885_), .C(decoded_rs1_2_bF_buf5_), .Y(_9889_) );
OAI21X1 OAI21X1_2089 ( .A(_7391_), .B(decoded_rs1_0_bF_buf55_), .C(_7556__bF_buf40), .Y(_9890_) );
AOI21X1 AOI21X1_675 ( .A(cpuregs_25_[29]), .B(decoded_rs1_0_bF_buf54_), .C(_9890_), .Y(_9891_) );
INVX1 INVX1_834 ( .A(cpuregs_27_[29]), .Y(_9892_) );
OAI21X1 OAI21X1_2090 ( .A(_9892_), .B(_7569__bF_buf30), .C(decoded_rs1_1_bF_buf33_), .Y(_9893_) );
AOI21X1 AOI21X1_676 ( .A(cpuregs_26_[29]), .B(_7569__bF_buf29), .C(_9893_), .Y(_9894_) );
OAI21X1 OAI21X1_2091 ( .A(_9894_), .B(_9891_), .C(_7560__bF_buf12), .Y(_9895_) );
AOI21X1 AOI21X1_677 ( .A(_9889_), .B(_9895_), .C(_7561__bF_buf1), .Y(_9896_) );
OAI21X1 OAI21X1_2092 ( .A(_9883_), .B(_9896_), .C(decoded_rs1_4_bF_buf4_), .Y(_9897_) );
NOR2X1 NOR2X1_872 ( .A(_7379_), .B(_7569__bF_buf28), .Y(_9898_) );
INVX1 INVX1_835 ( .A(cpuregs_8_[29]), .Y(_9899_) );
OAI21X1 OAI21X1_2093 ( .A(_9899_), .B(decoded_rs1_0_bF_buf53_), .C(_7556__bF_buf39), .Y(_9900_) );
AND2X2 AND2X2_148 ( .A(_7569__bF_buf27), .B(cpuregs_10_[29]), .Y(_9901_) );
INVX1 INVX1_836 ( .A(cpuregs_11_[29]), .Y(_9902_) );
OAI21X1 OAI21X1_2094 ( .A(_9902_), .B(_7569__bF_buf26), .C(decoded_rs1_1_bF_buf32_), .Y(_9903_) );
OAI22X1 OAI22X1_209 ( .A(_9900_), .B(_9898_), .C(_9903_), .D(_9901_), .Y(_9904_) );
NOR2X1 NOR2X1_873 ( .A(decoded_rs1_2_bF_buf4_), .B(_9904_), .Y(_9905_) );
NOR2X1 NOR2X1_874 ( .A(_7372_), .B(_7569__bF_buf25), .Y(_9906_) );
INVX1 INVX1_837 ( .A(cpuregs_12_[29]), .Y(_9907_) );
OAI21X1 OAI21X1_2095 ( .A(_9907_), .B(decoded_rs1_0_bF_buf52_), .C(_7556__bF_buf38), .Y(_9908_) );
AND2X2 AND2X2_149 ( .A(_7569__bF_buf24), .B(cpuregs_14_[29]), .Y(_9909_) );
INVX1 INVX1_838 ( .A(cpuregs_15_[29]), .Y(_9910_) );
OAI21X1 OAI21X1_2096 ( .A(_9910_), .B(_7569__bF_buf23), .C(decoded_rs1_1_bF_buf31_), .Y(_9911_) );
OAI22X1 OAI22X1_210 ( .A(_9908_), .B(_9906_), .C(_9911_), .D(_9909_), .Y(_9912_) );
OAI21X1 OAI21X1_2097 ( .A(_9912_), .B(_7560__bF_buf11), .C(decoded_rs1_3_bF_buf3_), .Y(_9913_) );
INVX1 INVX1_839 ( .A(cpuregs_4_[29]), .Y(_9914_) );
NAND2X1 NAND2X1_602 ( .A(cpuregs_6_[29]), .B(decoded_rs1_1_bF_buf30_), .Y(_9915_) );
OAI21X1 OAI21X1_2098 ( .A(_9914_), .B(decoded_rs1_1_bF_buf29_), .C(_9915_), .Y(_9916_) );
MUX2X1 MUX2X1_197 ( .A(cpuregs_7_[29]), .B(cpuregs_5_[29]), .S(decoded_rs1_1_bF_buf28_), .Y(_9917_) );
OAI21X1 OAI21X1_2099 ( .A(_9917_), .B(_7569__bF_buf22), .C(decoded_rs1_2_bF_buf3_), .Y(_9918_) );
AOI21X1 AOI21X1_678 ( .A(_7569__bF_buf21), .B(_9916_), .C(_9918_), .Y(_9919_) );
INVX1 INVX1_840 ( .A(cpuregs_0_[29]), .Y(_9920_) );
NAND2X1 NAND2X1_603 ( .A(cpuregs_2_[29]), .B(decoded_rs1_1_bF_buf27_), .Y(_9921_) );
OAI21X1 OAI21X1_2100 ( .A(_9920_), .B(decoded_rs1_1_bF_buf26_), .C(_9921_), .Y(_9922_) );
MUX2X1 MUX2X1_198 ( .A(cpuregs_3_[29]), .B(cpuregs_1_[29]), .S(decoded_rs1_1_bF_buf25_), .Y(_9923_) );
OAI21X1 OAI21X1_2101 ( .A(_9923_), .B(_7569__bF_buf20), .C(_7560__bF_buf10), .Y(_9924_) );
AOI21X1 AOI21X1_679 ( .A(_7569__bF_buf19), .B(_9922_), .C(_9924_), .Y(_9925_) );
OAI21X1 OAI21X1_2102 ( .A(_9919_), .B(_9925_), .C(_7561__bF_buf0), .Y(_9926_) );
OAI21X1 OAI21X1_2103 ( .A(_9905_), .B(_9913_), .C(_9926_), .Y(_9927_) );
AOI21X1 AOI21X1_680 ( .A(_7552__bF_buf3), .B(_9927_), .C(_7586__bF_buf2), .Y(_9928_) );
AOI22X1 AOI22X1_101 ( .A(reg_pc_29_), .B(_7551__bF_buf0), .C(_9928_), .D(_9897_), .Y(_9929_) );
NOR2X1 NOR2X1_875 ( .A(_4538__bF_buf2), .B(_9929_), .Y(_9930_) );
NOR2X1 NOR2X1_876 ( .A(_5027_), .B(_7700__bF_buf1), .Y(_9931_) );
AOI21X1 AOI21X1_681 ( .A(_10734__28_), .B(_8139_), .C(_4580__bF_buf2), .Y(_9932_) );
OAI21X1 OAI21X1_2104 ( .A(_4998_), .B(_7698__bF_buf2), .C(_9932_), .Y(_9933_) );
OAI21X1 OAI21X1_2105 ( .A(_9931_), .B(_9849_), .C(_9933_), .Y(_9934_) );
OAI21X1 OAI21X1_2106 ( .A(_7627_), .B(_5009_), .C(resetn_bF_buf5), .Y(_9935_) );
AOI21X1 AOI21X1_682 ( .A(_10734__29_), .B(_4597__bF_buf2), .C(_9935_), .Y(_9936_) );
OAI21X1 OAI21X1_2107 ( .A(_7697__bF_buf1), .B(_9934_), .C(_9936_), .Y(_9937_) );
OR2X2 OR2X2_21 ( .A(_9930_), .B(_9937_), .Y(_9938_) );
AOI21X1 AOI21X1_683 ( .A(_9869_), .B(_9868_), .C(_9938_), .Y(_9939_) );
AOI22X1 AOI22X1_102 ( .A(_4426__bF_buf2), .B(_5009_), .C(_9939_), .D(_9867_), .Y(_81__29_) );
NAND2X1 NAND2X1_604 ( .A(_9772_), .B(_9861_), .Y(_9940_) );
AOI21X1 AOI21X1_684 ( .A(_9771_), .B(_9861_), .C(_9860_), .Y(_9941_) );
OAI21X1 OAI21X1_2108 ( .A(_9775_), .B(_9940_), .C(_9941_), .Y(_9942_) );
INVX1 INVX1_841 ( .A(decoded_imm_30_), .Y(_9943_) );
NAND2X1 NAND2X1_605 ( .A(_4998_), .B(_9943_), .Y(_9944_) );
NOR2X1 NOR2X1_877 ( .A(_4998_), .B(_9943_), .Y(_9945_) );
INVX1 INVX1_842 ( .A(_9945_), .Y(_9946_) );
AND2X2 AND2X2_150 ( .A(_9946_), .B(_9944_), .Y(_9947_) );
NOR2X1 NOR2X1_878 ( .A(_9947_), .B(_9942_), .Y(_9948_) );
INVX1 INVX1_843 ( .A(_9940_), .Y(_9949_) );
OAI21X1 OAI21X1_2109 ( .A(_9766_), .B(_9768_), .C(_9949_), .Y(_9950_) );
INVX1 INVX1_844 ( .A(_9947_), .Y(_9951_) );
AOI21X1 AOI21X1_685 ( .A(_9941_), .B(_9950_), .C(_9951_), .Y(_9952_) );
OAI21X1 OAI21X1_2110 ( .A(_9948_), .B(_9952_), .C(_7624__bF_buf4), .Y(_9953_) );
AOI21X1 AOI21X1_686 ( .A(_4998_), .B(_7623__bF_buf0), .C(_4587__bF_buf1), .Y(_9954_) );
NAND2X1 NAND2X1_606 ( .A(_9954_), .B(_9953_), .Y(_9955_) );
OAI21X1 OAI21X1_2111 ( .A(_9948_), .B(_9952_), .C(_7632__bF_buf3), .Y(_9956_) );
AOI21X1 AOI21X1_687 ( .A(_4998_), .B(_7631__bF_buf1), .C(_7629__bF_buf3), .Y(_9957_) );
AND2X2 AND2X2_151 ( .A(cpuregs_1_[30]), .B(decoded_rs1_0_bF_buf51_), .Y(_9958_) );
INVX1 INVX1_845 ( .A(cpuregs_0_[30]), .Y(_9959_) );
OAI21X1 OAI21X1_2112 ( .A(_9959_), .B(decoded_rs1_0_bF_buf50_), .C(_7556__bF_buf37), .Y(_9960_) );
NOR2X1 NOR2X1_879 ( .A(decoded_rs1_0_bF_buf49_), .B(_7443_), .Y(_9961_) );
INVX1 INVX1_846 ( .A(cpuregs_3_[30]), .Y(_9962_) );
OAI21X1 OAI21X1_2113 ( .A(_9962_), .B(_7569__bF_buf18), .C(decoded_rs1_1_bF_buf24_), .Y(_9963_) );
OAI22X1 OAI22X1_211 ( .A(_9960_), .B(_9958_), .C(_9963_), .D(_9961_), .Y(_9964_) );
NOR2X1 NOR2X1_880 ( .A(decoded_rs1_2_bF_buf2_), .B(_9964_), .Y(_9965_) );
AND2X2 AND2X2_152 ( .A(cpuregs_5_[30]), .B(decoded_rs1_0_bF_buf48_), .Y(_9966_) );
INVX1 INVX1_847 ( .A(cpuregs_4_[30]), .Y(_9967_) );
OAI21X1 OAI21X1_2114 ( .A(_9967_), .B(decoded_rs1_0_bF_buf47_), .C(_7556__bF_buf36), .Y(_9968_) );
NOR2X1 NOR2X1_881 ( .A(decoded_rs1_0_bF_buf46_), .B(_7437_), .Y(_9969_) );
INVX1 INVX1_848 ( .A(cpuregs_7_[30]), .Y(_9970_) );
OAI21X1 OAI21X1_2115 ( .A(_9970_), .B(_7569__bF_buf17), .C(decoded_rs1_1_bF_buf23_), .Y(_9971_) );
OAI22X1 OAI22X1_212 ( .A(_9968_), .B(_9966_), .C(_9971_), .D(_9969_), .Y(_9972_) );
OAI21X1 OAI21X1_2116 ( .A(_9972_), .B(_7560__bF_buf9), .C(_7561__bF_buf6), .Y(_9973_) );
NOR2X1 NOR2X1_882 ( .A(_9965_), .B(_9973_), .Y(_9974_) );
NOR2X1 NOR2X1_883 ( .A(cpuregs_14_[30]), .B(_7556__bF_buf35), .Y(_9975_) );
OAI21X1 OAI21X1_2117 ( .A(cpuregs_12_[30]), .B(decoded_rs1_1_bF_buf22_), .C(_7569__bF_buf16), .Y(_9976_) );
NOR2X1 NOR2X1_884 ( .A(cpuregs_15_[30]), .B(_7556__bF_buf34), .Y(_9977_) );
OAI21X1 OAI21X1_2118 ( .A(cpuregs_13_[30]), .B(decoded_rs1_1_bF_buf21_), .C(decoded_rs1_0_bF_buf45_), .Y(_9978_) );
OAI22X1 OAI22X1_213 ( .A(_9975_), .B(_9976_), .C(_9977_), .D(_9978_), .Y(_9979_) );
NOR2X1 NOR2X1_885 ( .A(cpuregs_10_[30]), .B(_7556__bF_buf33), .Y(_9980_) );
OAI21X1 OAI21X1_2119 ( .A(cpuregs_8_[30]), .B(decoded_rs1_1_bF_buf20_), .C(_7569__bF_buf15), .Y(_9981_) );
NOR2X1 NOR2X1_886 ( .A(cpuregs_11_[30]), .B(_7556__bF_buf32), .Y(_9982_) );
OAI21X1 OAI21X1_2120 ( .A(cpuregs_9_[30]), .B(decoded_rs1_1_bF_buf19_), .C(decoded_rs1_0_bF_buf44_), .Y(_9983_) );
OAI22X1 OAI22X1_214 ( .A(_9980_), .B(_9981_), .C(_9982_), .D(_9983_), .Y(_9984_) );
MUX2X1 MUX2X1_199 ( .A(_9984_), .B(_9979_), .S(_7560__bF_buf8), .Y(_9985_) );
AND2X2 AND2X2_153 ( .A(_9985_), .B(decoded_rs1_3_bF_buf2_), .Y(_9986_) );
OAI21X1 OAI21X1_2121 ( .A(_9986_), .B(_9974_), .C(_7552__bF_buf2), .Y(_9987_) );
AOI21X1 AOI21X1_688 ( .A(_7455_), .B(_7556__bF_buf31), .C(decoded_rs1_0_bF_buf43_), .Y(_9988_) );
OAI21X1 OAI21X1_2122 ( .A(cpuregs_30_[30]), .B(_7556__bF_buf30), .C(_9988_), .Y(_9989_) );
AOI21X1 AOI21X1_689 ( .A(_7452_), .B(_7556__bF_buf29), .C(_7569__bF_buf14), .Y(_9990_) );
OAI21X1 OAI21X1_2123 ( .A(cpuregs_31_[30]), .B(_7556__bF_buf28), .C(_9990_), .Y(_9991_) );
AOI21X1 AOI21X1_690 ( .A(_9989_), .B(_9991_), .C(_7560__bF_buf7), .Y(_9992_) );
AND2X2 AND2X2_154 ( .A(cpuregs_17_[30]), .B(decoded_rs1_0_bF_buf42_), .Y(_9993_) );
INVX1 INVX1_849 ( .A(cpuregs_16_[30]), .Y(_9994_) );
OAI21X1 OAI21X1_2124 ( .A(_9994_), .B(decoded_rs1_0_bF_buf41_), .C(_7556__bF_buf27), .Y(_9995_) );
AND2X2 AND2X2_155 ( .A(_7569__bF_buf13), .B(cpuregs_18_[30]), .Y(_9996_) );
INVX1 INVX1_850 ( .A(cpuregs_19_[30]), .Y(_9997_) );
OAI21X1 OAI21X1_2125 ( .A(_9997_), .B(_7569__bF_buf12), .C(decoded_rs1_1_bF_buf18_), .Y(_9998_) );
OAI22X1 OAI22X1_215 ( .A(_9995_), .B(_9993_), .C(_9998_), .D(_9996_), .Y(_9999_) );
NOR2X1 NOR2X1_887 ( .A(decoded_rs1_2_bF_buf1_), .B(_9999_), .Y(_10000_) );
NOR2X1 NOR2X1_888 ( .A(_7425_), .B(_7569__bF_buf11), .Y(_10001_) );
OAI21X1 OAI21X1_2126 ( .A(_7422_), .B(decoded_rs1_0_bF_buf40_), .C(_7556__bF_buf26), .Y(_10002_) );
NOR2X1 NOR2X1_889 ( .A(decoded_rs1_0_bF_buf39_), .B(_7429_), .Y(_10003_) );
OAI21X1 OAI21X1_2127 ( .A(_7432_), .B(_7569__bF_buf10), .C(decoded_rs1_1_bF_buf17_), .Y(_10004_) );
OAI22X1 OAI22X1_216 ( .A(_10002_), .B(_10001_), .C(_10004_), .D(_10003_), .Y(_10005_) );
OAI21X1 OAI21X1_2128 ( .A(_10005_), .B(_7560__bF_buf6), .C(_7561__bF_buf5), .Y(_10006_) );
AND2X2 AND2X2_156 ( .A(cpuregs_25_[30]), .B(decoded_rs1_0_bF_buf38_), .Y(_10007_) );
OAI21X1 OAI21X1_2129 ( .A(_7460_), .B(decoded_rs1_0_bF_buf37_), .C(_7556__bF_buf25), .Y(_10008_) );
AND2X2 AND2X2_157 ( .A(_7569__bF_buf9), .B(cpuregs_26_[30]), .Y(_10009_) );
OAI21X1 OAI21X1_2130 ( .A(_7463_), .B(_7569__bF_buf8), .C(decoded_rs1_1_bF_buf16_), .Y(_10010_) );
OAI22X1 OAI22X1_217 ( .A(_10008_), .B(_10007_), .C(_10010_), .D(_10009_), .Y(_10011_) );
OAI21X1 OAI21X1_2131 ( .A(_10011_), .B(decoded_rs1_2_bF_buf0_), .C(decoded_rs1_3_bF_buf1_), .Y(_10012_) );
OAI22X1 OAI22X1_218 ( .A(_10006_), .B(_10000_), .C(_9992_), .D(_10012_), .Y(_10013_) );
AOI21X1 AOI21X1_691 ( .A(decoded_rs1_4_bF_buf3_), .B(_10013_), .C(_7586__bF_buf1), .Y(_10014_) );
AOI22X1 AOI22X1_103 ( .A(reg_pc_30_), .B(_7551__bF_buf3), .C(_10014_), .D(_9987_), .Y(_10015_) );
NOR2X1 NOR2X1_890 ( .A(_4538__bF_buf1), .B(_10015_), .Y(_10016_) );
INVX1 INVX1_851 ( .A(_9755_), .Y(_10017_) );
AOI21X1 AOI21X1_692 ( .A(_10734__29_), .B(_8139_), .C(_4580__bF_buf1), .Y(_10018_) );
OAI21X1 OAI21X1_2132 ( .A(_4991_), .B(_7698__bF_buf1), .C(_10018_), .Y(_10019_) );
OAI21X1 OAI21X1_2133 ( .A(_10017_), .B(_9849_), .C(_10019_), .Y(_10020_) );
OAI21X1 OAI21X1_2134 ( .A(_7627_), .B(_4998_), .C(resetn_bF_buf4), .Y(_10021_) );
AOI21X1 AOI21X1_693 ( .A(_10734__30_), .B(_4597__bF_buf1), .C(_10021_), .Y(_10022_) );
OAI21X1 OAI21X1_2135 ( .A(_7697__bF_buf0), .B(_10020_), .C(_10022_), .Y(_10023_) );
OR2X2 OR2X2_22 ( .A(_10023_), .B(_10016_), .Y(_10024_) );
AOI21X1 AOI21X1_694 ( .A(_9957_), .B(_9956_), .C(_10024_), .Y(_10025_) );
AOI22X1 AOI22X1_104 ( .A(_4426__bF_buf1), .B(_4998_), .C(_10025_), .D(_9955_), .Y(_81__30_) );
NAND2X1 NAND2X1_607 ( .A(_9947_), .B(_9942_), .Y(_10026_) );
XNOR2X1 XNOR2X1_14 ( .A(_10734__31_), .B(decoded_imm_31_), .Y(_10027_) );
INVX1 INVX1_852 ( .A(_10027_), .Y(_10028_) );
NAND3X1 NAND3X1_54 ( .A(_9946_), .B(_10028_), .C(_10026_), .Y(_10029_) );
OAI21X1 OAI21X1_2136 ( .A(_9952_), .B(_9945_), .C(_10027_), .Y(_10030_) );
NAND2X1 NAND2X1_608 ( .A(_10030_), .B(_10029_), .Y(_10031_) );
AOI21X1 AOI21X1_695 ( .A(_4991_), .B(_7623__bF_buf4), .C(_4587__bF_buf0), .Y(_10032_) );
OAI21X1 OAI21X1_2137 ( .A(_10031_), .B(_7623__bF_buf3), .C(_10032_), .Y(_10033_) );
NAND3X1 NAND3X1_55 ( .A(_7632__bF_buf2), .B(_10030_), .C(_10029_), .Y(_10034_) );
AOI21X1 AOI21X1_696 ( .A(_4991_), .B(_7631__bF_buf0), .C(_7629__bF_buf2), .Y(_10035_) );
NOR2X1 NOR2X1_891 ( .A(cpuregs_4_[31]), .B(decoded_rs1_0_bF_buf36_), .Y(_10036_) );
OAI21X1 OAI21X1_2138 ( .A(_7569__bF_buf7), .B(cpuregs_5_[31]), .C(_7556__bF_buf24), .Y(_10037_) );
NOR2X1 NOR2X1_892 ( .A(cpuregs_7_[31]), .B(_7569__bF_buf6), .Y(_10038_) );
OAI21X1 OAI21X1_2139 ( .A(cpuregs_6_[31]), .B(decoded_rs1_0_bF_buf35_), .C(decoded_rs1_1_bF_buf15_), .Y(_10039_) );
OAI22X1 OAI22X1_219 ( .A(_10038_), .B(_10039_), .C(_10037_), .D(_10036_), .Y(_10040_) );
NAND2X1 NAND2X1_609 ( .A(decoded_rs1_2_bF_buf12_), .B(_10040_), .Y(_10041_) );
OAI21X1 OAI21X1_2140 ( .A(_7569__bF_buf5), .B(cpuregs_1_[31]), .C(_7556__bF_buf23), .Y(_10042_) );
AOI21X1 AOI21X1_697 ( .A(_7484_), .B(_7569__bF_buf4), .C(_10042_), .Y(_10043_) );
INVX1 INVX1_853 ( .A(cpuregs_3_[31]), .Y(_10044_) );
OAI21X1 OAI21X1_2141 ( .A(cpuregs_2_[31]), .B(decoded_rs1_0_bF_buf34_), .C(decoded_rs1_1_bF_buf14_), .Y(_10045_) );
AOI21X1 AOI21X1_698 ( .A(_10044_), .B(decoded_rs1_0_bF_buf33_), .C(_10045_), .Y(_10046_) );
OAI21X1 OAI21X1_2142 ( .A(_10043_), .B(_10046_), .C(_7560__bF_buf5), .Y(_10047_) );
AOI21X1 AOI21X1_699 ( .A(_10041_), .B(_10047_), .C(decoded_rs1_3_bF_buf0_), .Y(_10048_) );
OAI21X1 OAI21X1_2143 ( .A(_7508_), .B(decoded_rs1_0_bF_buf32_), .C(decoded_rs1_1_bF_buf13_), .Y(_10049_) );
AOI21X1 AOI21X1_700 ( .A(cpuregs_15_[31]), .B(decoded_rs1_0_bF_buf31_), .C(_10049_), .Y(_10050_) );
NOR2X1 NOR2X1_893 ( .A(decoded_rs1_0_bF_buf30_), .B(_7510_), .Y(_10051_) );
OAI21X1 OAI21X1_2144 ( .A(_7505_), .B(_7569__bF_buf3), .C(_7556__bF_buf22), .Y(_10052_) );
OAI21X1 OAI21X1_2145 ( .A(_10052_), .B(_10051_), .C(decoded_rs1_2_bF_buf11_), .Y(_10053_) );
AOI21X1 AOI21X1_701 ( .A(cpuregs_10_[31]), .B(_7569__bF_buf2), .C(_7556__bF_buf21), .Y(_10054_) );
OAI21X1 OAI21X1_2146 ( .A(_7501_), .B(_7569__bF_buf1), .C(_10054_), .Y(_10055_) );
AOI21X1 AOI21X1_702 ( .A(cpuregs_8_[31]), .B(_7569__bF_buf0), .C(decoded_rs1_1_bF_buf12_), .Y(_10056_) );
OAI21X1 OAI21X1_2147 ( .A(_7498_), .B(_7569__bF_buf48), .C(_10056_), .Y(_10057_) );
NAND3X1 NAND3X1_56 ( .A(_7560__bF_buf4), .B(_10055_), .C(_10057_), .Y(_10058_) );
OAI21X1 OAI21X1_2148 ( .A(_10050_), .B(_10053_), .C(_10058_), .Y(_10059_) );
AOI21X1 AOI21X1_703 ( .A(decoded_rs1_3_bF_buf6_), .B(_10059_), .C(_10048_), .Y(_10060_) );
AND2X2 AND2X2_158 ( .A(_10060_), .B(_7552__bF_buf1), .Y(_10061_) );
NOR2X1 NOR2X1_894 ( .A(cpuregs_16_[31]), .B(decoded_rs1_0_bF_buf29_), .Y(_10062_) );
OAI21X1 OAI21X1_2149 ( .A(_7569__bF_buf47), .B(cpuregs_17_[31]), .C(_7556__bF_buf20), .Y(_10063_) );
NOR2X1 NOR2X1_895 ( .A(cpuregs_19_[31]), .B(_7569__bF_buf46), .Y(_10064_) );
OAI21X1 OAI21X1_2150 ( .A(cpuregs_18_[31]), .B(decoded_rs1_0_bF_buf28_), .C(decoded_rs1_1_bF_buf11_), .Y(_10065_) );
OAI22X1 OAI22X1_220 ( .A(_10064_), .B(_10065_), .C(_10063_), .D(_10062_), .Y(_10066_) );
NOR2X1 NOR2X1_896 ( .A(decoded_rs1_2_bF_buf10_), .B(_10066_), .Y(_10067_) );
NOR2X1 NOR2X1_897 ( .A(cpuregs_20_[31]), .B(decoded_rs1_0_bF_buf27_), .Y(_10068_) );
OAI21X1 OAI21X1_2151 ( .A(_7569__bF_buf45), .B(cpuregs_21_[31]), .C(_7556__bF_buf19), .Y(_10069_) );
NOR2X1 NOR2X1_898 ( .A(cpuregs_23_[31]), .B(_7569__bF_buf44), .Y(_10070_) );
OAI21X1 OAI21X1_2152 ( .A(cpuregs_22_[31]), .B(decoded_rs1_0_bF_buf26_), .C(decoded_rs1_1_bF_buf10_), .Y(_10071_) );
OAI22X1 OAI22X1_221 ( .A(_10070_), .B(_10071_), .C(_10069_), .D(_10068_), .Y(_10072_) );
OAI21X1 OAI21X1_2153 ( .A(_10072_), .B(_7560__bF_buf3), .C(_7561__bF_buf4), .Y(_10073_) );
NAND2X1 NAND2X1_610 ( .A(cpuregs_29_[31]), .B(decoded_rs1_0_bF_buf25_), .Y(_10074_) );
OAI21X1 OAI21X1_2154 ( .A(_7538_), .B(decoded_rs1_0_bF_buf24_), .C(_10074_), .Y(_10075_) );
NAND2X1 NAND2X1_611 ( .A(cpuregs_31_[31]), .B(decoded_rs1_0_bF_buf23_), .Y(_10076_) );
OAI21X1 OAI21X1_2155 ( .A(_7541_), .B(decoded_rs1_0_bF_buf22_), .C(_10076_), .Y(_10077_) );
MUX2X1 MUX2X1_200 ( .A(_10077_), .B(_10075_), .S(decoded_rs1_1_bF_buf9_), .Y(_10078_) );
NOR2X1 NOR2X1_899 ( .A(_7560__bF_buf2), .B(_10078_), .Y(_10079_) );
OAI21X1 OAI21X1_2156 ( .A(_7531_), .B(decoded_rs1_0_bF_buf21_), .C(decoded_rs1_1_bF_buf8_), .Y(_10080_) );
AOI21X1 AOI21X1_704 ( .A(cpuregs_27_[31]), .B(decoded_rs1_0_bF_buf20_), .C(_10080_), .Y(_10081_) );
AND2X2 AND2X2_159 ( .A(cpuregs_25_[31]), .B(decoded_rs1_0_bF_buf19_), .Y(_10082_) );
OAI21X1 OAI21X1_2157 ( .A(_7535_), .B(decoded_rs1_0_bF_buf18_), .C(_7556__bF_buf18), .Y(_10083_) );
OAI21X1 OAI21X1_2158 ( .A(_10083_), .B(_10082_), .C(_7560__bF_buf1), .Y(_10084_) );
NOR2X1 NOR2X1_900 ( .A(_10081_), .B(_10084_), .Y(_10085_) );
OAI21X1 OAI21X1_2159 ( .A(_10079_), .B(_10085_), .C(decoded_rs1_3_bF_buf5_), .Y(_10086_) );
OAI21X1 OAI21X1_2160 ( .A(_10067_), .B(_10073_), .C(_10086_), .Y(_10087_) );
OAI21X1 OAI21X1_2161 ( .A(_10087_), .B(_7552__bF_buf0), .C(_7587_), .Y(_10088_) );
OAI22X1 OAI22X1_222 ( .A(_4907_), .B(_7643_), .C(_10061_), .D(_10088_), .Y(_10089_) );
NAND2X1 NAND2X1_612 ( .A(cpu_state_2_bF_buf3_), .B(_10089_), .Y(_10090_) );
OAI21X1 OAI21X1_2162 ( .A(_4597__bF_buf0), .B(_8855_), .C(_10734__31_), .Y(_10091_) );
OAI21X1 OAI21X1_2163 ( .A(_4998_), .B(_7700__bF_buf0), .C(_4579__bF_buf3), .Y(_10092_) );
OAI21X1 OAI21X1_2164 ( .A(_4578_), .B(reg_sh_4_), .C(_9850_), .Y(_10093_) );
NAND2X1 NAND2X1_613 ( .A(_10093_), .B(_10092_), .Y(_10094_) );
NAND2X1 NAND2X1_614 ( .A(_9848_), .B(_10094_), .Y(_10095_) );
AOI21X1 AOI21X1_705 ( .A(_10095_), .B(_4584_), .C(_4426__bF_buf0), .Y(_10096_) );
NAND3X1 NAND3X1_57 ( .A(_10091_), .B(_10096_), .C(_10090_), .Y(_10097_) );
AOI21X1 AOI21X1_706 ( .A(_10035_), .B(_10034_), .C(_10097_), .Y(_10098_) );
AOI22X1 AOI22X1_105 ( .A(_4426__bF_buf11), .B(_4991_), .C(_10098_), .D(_10033_), .Y(_81__31_) );
NOR2X1 NOR2X1_901 ( .A(_4431__bF_buf4), .B(_4605__bF_buf4), .Y(_10099_) );
INVX1 INVX1_854 ( .A(decoded_imm_uj_0_), .Y(_10100_) );
NOR2X1 NOR2X1_902 ( .A(_4499__bF_buf4), .B(_10100_), .Y(_10101_) );
NAND2X1 NAND2X1_615 ( .A(_10099__bF_buf3), .B(_10101_), .Y(_10102_) );
NAND2X1 NAND2X1_616 ( .A(latched_branch), .B(latched_store), .Y(_10103_) );
OAI21X1 OAI21X1_2165 ( .A(_10103__bF_buf6), .B(_4431__bF_buf3), .C(reg_next_pc_0_), .Y(_10104_) );
OAI21X1 OAI21X1_2166 ( .A(_10102_), .B(_10104_), .C(resetn_bF_buf3), .Y(_10105_) );
AOI21X1 AOI21X1_707 ( .A(_10102_), .B(_10104_), .C(_10105_), .Y(_80__0_) );
NAND2X1 NAND2X1_617 ( .A(reg_next_pc_1_), .B(_4431__bF_buf2), .Y(_10106_) );
NOR2X1 NOR2X1_903 ( .A(_4499__bF_buf3), .B(_4605__bF_buf3), .Y(_10107_) );
INVX1 INVX1_855 ( .A(_10107_), .Y(_10108_) );
INVX1 INVX1_856 ( .A(latched_branch), .Y(_10109_) );
OAI21X1 OAI21X1_2167 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_0_), .Y(_10110_) );
NOR2X1 NOR2X1_904 ( .A(_10100_), .B(_10110_), .Y(_10111_) );
INVX1 INVX1_857 ( .A(decoded_imm_uj_1_), .Y(_10112_) );
AOI21X1 AOI21X1_708 ( .A(latched_branch), .B(latched_store), .C(reg_next_pc_1_), .Y(_10113_) );
INVX1 INVX1_858 ( .A(_10113_), .Y(_10114_) );
OAI21X1 OAI21X1_2168 ( .A(_4932_), .B(_10103__bF_buf5), .C(_10114_), .Y(_10115_) );
NAND2X1 NAND2X1_618 ( .A(_10112_), .B(_10115_), .Y(_10116_) );
MUX2X1 MUX2X1_201 ( .A(alu_out_q_1_), .B(reg_out_1_), .S(latched_stalu_bF_buf0), .Y(_10117_) );
AND2X2 AND2X2_160 ( .A(latched_branch), .B(latched_store), .Y(_10118_) );
AOI21X1 AOI21X1_709 ( .A(_10118__bF_buf4), .B(_10117_), .C(_10113_), .Y(_10119_) );
NAND2X1 NAND2X1_619 ( .A(decoded_imm_uj_1_), .B(_10119_), .Y(_10120_) );
NAND2X1 NAND2X1_620 ( .A(_10120_), .B(_10116_), .Y(_10121_) );
XNOR2X1 XNOR2X1_15 ( .A(_10121_), .B(_10111_), .Y(_10122_) );
INVX1 INVX1_859 ( .A(_10099__bF_buf2), .Y(_10123_) );
NAND2X1 NAND2X1_621 ( .A(cpu_state_1_bF_buf0_), .B(_10119_), .Y(_10124_) );
OAI21X1 OAI21X1_2169 ( .A(_4499__bF_buf2), .B(_10123__bF_buf4), .C(_10124_), .Y(_10125_) );
OAI21X1 OAI21X1_2170 ( .A(_10122_), .B(_10108_), .C(_10125_), .Y(_10126_) );
AOI21X1 AOI21X1_710 ( .A(_10106_), .B(_10126_), .C(_4426__bF_buf10), .Y(_80__1_) );
AND2X2 AND2X2_161 ( .A(_10119_), .B(decoded_imm_uj_1_), .Y(_10127_) );
AOI21X1 AOI21X1_711 ( .A(_10111_), .B(_10116_), .C(_10127_), .Y(_10128_) );
MUX2X1 MUX2X1_202 ( .A(alu_out_q_2_), .B(reg_out_2_), .S(latched_stalu_bF_buf6), .Y(_10129_) );
OAI21X1 OAI21X1_2171 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_2_), .Y(_10130_) );
OAI21X1 OAI21X1_2172 ( .A(_10129_), .B(_10103__bF_buf4), .C(_10130_), .Y(_10131_) );
NAND2X1 NAND2X1_622 ( .A(decoded_imm_uj_2_), .B(_10131_), .Y(_10132_) );
INVX1 INVX1_860 ( .A(decoded_imm_uj_2_), .Y(_10133_) );
MUX2X1 MUX2X1_203 ( .A(_4939_), .B(reg_next_pc_2_), .S(_10118__bF_buf3), .Y(_10134_) );
NAND2X1 NAND2X1_623 ( .A(_10133_), .B(_10134_), .Y(_10135_) );
NAND2X1 NAND2X1_624 ( .A(_10132_), .B(_10135_), .Y(_10136_) );
AOI21X1 AOI21X1_712 ( .A(_10136_), .B(_10128_), .C(_10108_), .Y(_10137_) );
OAI21X1 OAI21X1_2173 ( .A(_10128_), .B(_10136_), .C(_10137_), .Y(_10138_) );
OAI21X1 OAI21X1_2174 ( .A(_10134_), .B(decoder_trigger_bF_buf2), .C(cpu_state_1_bF_buf5_), .Y(_10139_) );
AOI21X1 AOI21X1_713 ( .A(_4606_), .B(_10134_), .C(_10139_), .Y(_10140_) );
OAI21X1 OAI21X1_2175 ( .A(cpu_state_1_bF_buf4_), .B(reg_next_pc_2_), .C(resetn_bF_buf2), .Y(_10141_) );
AOI21X1 AOI21X1_714 ( .A(_10140_), .B(_10138_), .C(_10141_), .Y(_80__2_) );
NAND2X1 NAND2X1_625 ( .A(reg_next_pc_3_), .B(_4431__bF_buf1), .Y(_10142_) );
MUX2X1 MUX2X1_204 ( .A(_4947_), .B(reg_next_pc_3_), .S(_10118__bF_buf2), .Y(_10143_) );
NOR2X1 NOR2X1_905 ( .A(_4431__bF_buf0), .B(_10143_), .Y(_10144_) );
OAI21X1 OAI21X1_2176 ( .A(_10128_), .B(_10136_), .C(_10132_), .Y(_10145_) );
MUX2X1 MUX2X1_205 ( .A(alu_out_q_3_), .B(reg_out_3_), .S(latched_stalu_bF_buf5), .Y(_10146_) );
OAI21X1 OAI21X1_2177 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_3_), .Y(_10147_) );
OAI21X1 OAI21X1_2178 ( .A(_10146_), .B(_10103__bF_buf3), .C(_10147_), .Y(_10148_) );
NOR2X1 NOR2X1_906 ( .A(decoded_imm_uj_3_), .B(_10148_), .Y(_10149_) );
INVX1 INVX1_861 ( .A(decoded_imm_uj_3_), .Y(_10150_) );
NOR2X1 NOR2X1_907 ( .A(_10150_), .B(_10143_), .Y(_10151_) );
NOR2X1 NOR2X1_908 ( .A(_10149_), .B(_10151_), .Y(_10152_) );
AOI21X1 AOI21X1_715 ( .A(_10152_), .B(_10145_), .C(_4499__bF_buf1), .Y(_10153_) );
OAI21X1 OAI21X1_2179 ( .A(_10145_), .B(_10152_), .C(_10153_), .Y(_10154_) );
NAND2X1 NAND2X1_626 ( .A(_10131_), .B(_10148_), .Y(_10155_) );
NAND2X1 NAND2X1_627 ( .A(_10134_), .B(_10143_), .Y(_10156_) );
AOI21X1 AOI21X1_716 ( .A(_10155_), .B(_10156_), .C(_4605__bF_buf2), .Y(_10157_) );
OAI21X1 OAI21X1_2180 ( .A(_10107_), .B(_10157_), .C(_10154_), .Y(_10158_) );
OAI21X1 OAI21X1_2181 ( .A(_10099__bF_buf1), .B(_10144_), .C(_10158_), .Y(_10159_) );
AOI21X1 AOI21X1_717 ( .A(_10142_), .B(_10159_), .C(_4426__bF_buf9), .Y(_80__3_) );
NAND2X1 NAND2X1_628 ( .A(reg_next_pc_4_), .B(_4431__bF_buf7), .Y(_10160_) );
MUX2X1 MUX2X1_206 ( .A(_4954_), .B(reg_next_pc_4_), .S(_10118__bF_buf1), .Y(_10161_) );
OAI21X1 OAI21X1_2182 ( .A(_10161_), .B(_4431__bF_buf6), .C(_10123__bF_buf3), .Y(_10162_) );
INVX1 INVX1_862 ( .A(decoded_imm_uj_4_), .Y(_10163_) );
MUX2X1 MUX2X1_207 ( .A(alu_out_q_4_), .B(reg_out_4_), .S(latched_stalu_bF_buf4), .Y(_10164_) );
OAI21X1 OAI21X1_2183 ( .A(_10109__bF_buf1), .B(_4639__bF_buf3), .C(reg_next_pc_4_), .Y(_10165_) );
OAI21X1 OAI21X1_2184 ( .A(_10164_), .B(_10103__bF_buf2), .C(_10165_), .Y(_10166_) );
XNOR2X1 XNOR2X1_16 ( .A(_10166_), .B(_10163_), .Y(_10167_) );
NAND2X1 NAND2X1_629 ( .A(decoded_imm_uj_3_), .B(_10148_), .Y(_10168_) );
OAI21X1 OAI21X1_2185 ( .A(_10149_), .B(_10132_), .C(_10168_), .Y(_10169_) );
INVX1 INVX1_863 ( .A(_10169_), .Y(_10170_) );
INVX1 INVX1_864 ( .A(_10111_), .Y(_10171_) );
NOR2X1 NOR2X1_909 ( .A(decoded_imm_uj_1_), .B(_10119_), .Y(_10172_) );
OAI21X1 OAI21X1_2186 ( .A(_10172_), .B(_10171_), .C(_10120_), .Y(_10173_) );
AND2X2 AND2X2_162 ( .A(_10135_), .B(_10132_), .Y(_10174_) );
NAND3X1 NAND3X1_58 ( .A(_10173_), .B(_10174_), .C(_10152_), .Y(_10175_) );
NAND2X1 NAND2X1_630 ( .A(_10170_), .B(_10175_), .Y(_10176_) );
OAI21X1 OAI21X1_2187 ( .A(_10176_), .B(_10167_), .C(instr_jal_bF_buf4), .Y(_10177_) );
AOI21X1 AOI21X1_718 ( .A(_10167_), .B(_10176_), .C(_10177_), .Y(_10178_) );
INVX1 INVX1_865 ( .A(_10155_), .Y(_10179_) );
NAND2X1 NAND2X1_631 ( .A(_10166_), .B(_10179_), .Y(_10180_) );
OAI21X1 OAI21X1_2188 ( .A(_10134_), .B(_10143_), .C(_10161_), .Y(_10181_) );
NAND2X1 NAND2X1_632 ( .A(_10181_), .B(_10180_), .Y(_10182_) );
OAI21X1 OAI21X1_2189 ( .A(_10182_), .B(instr_jal_bF_buf3), .C(decoder_trigger_bF_buf1), .Y(_10183_) );
OAI21X1 OAI21X1_2190 ( .A(_10178_), .B(_10183_), .C(_10162_), .Y(_10184_) );
AOI21X1 AOI21X1_719 ( .A(_10160_), .B(_10184_), .C(_4426__bF_buf8), .Y(_80__4_) );
NAND2X1 NAND2X1_633 ( .A(reg_next_pc_5_), .B(_4431__bF_buf5), .Y(_10185_) );
NAND2X1 NAND2X1_634 ( .A(decoded_imm_uj_4_), .B(_10166_), .Y(_10186_) );
XNOR2X1 XNOR2X1_17 ( .A(_10166_), .B(decoded_imm_uj_4_), .Y(_10187_) );
INVX1 INVX1_866 ( .A(_10176_), .Y(_10188_) );
OAI21X1 OAI21X1_2191 ( .A(_10188_), .B(_10187_), .C(_10186_), .Y(_10189_) );
INVX1 INVX1_867 ( .A(decoded_imm_uj_5_), .Y(_10190_) );
OAI21X1 OAI21X1_2192 ( .A(_10109__bF_buf0), .B(_4639__bF_buf2), .C(reg_next_pc_5_), .Y(_10191_) );
OAI21X1 OAI21X1_2193 ( .A(_4652_), .B(_10103__bF_buf1), .C(_10191_), .Y(_10192_) );
XNOR2X1 XNOR2X1_18 ( .A(_10192_), .B(_10190_), .Y(_10193_) );
OAI21X1 OAI21X1_2194 ( .A(_10189_), .B(_10193_), .C(instr_jal_bF_buf2), .Y(_10194_) );
AOI21X1 AOI21X1_720 ( .A(_10189_), .B(_10193_), .C(_10194_), .Y(_10195_) );
INVX1 INVX1_868 ( .A(_10192_), .Y(_10196_) );
NOR2X1 NOR2X1_910 ( .A(_10161_), .B(_10196_), .Y(_10197_) );
NAND2X1 NAND2X1_635 ( .A(_10179_), .B(_10197_), .Y(_10198_) );
OAI21X1 OAI21X1_2195 ( .A(_10155_), .B(_10161_), .C(_10196_), .Y(_10199_) );
NAND2X1 NAND2X1_636 ( .A(_10199_), .B(_10198_), .Y(_10200_) );
OAI21X1 OAI21X1_2196 ( .A(_10200_), .B(instr_jal_bF_buf1), .C(decoder_trigger_bF_buf0), .Y(_10201_) );
OAI21X1 OAI21X1_2197 ( .A(_10196_), .B(_4431__bF_buf4), .C(_10123__bF_buf2), .Y(_10202_) );
OAI21X1 OAI21X1_2198 ( .A(_10195_), .B(_10201_), .C(_10202_), .Y(_10203_) );
AOI21X1 AOI21X1_721 ( .A(_10185_), .B(_10203_), .C(_4426__bF_buf7), .Y(_80__5_) );
NAND2X1 NAND2X1_637 ( .A(reg_next_pc_6_), .B(_4431__bF_buf3), .Y(_10204_) );
OAI21X1 OAI21X1_2199 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_6_), .Y(_10205_) );
OAI21X1 OAI21X1_2200 ( .A(_4662_), .B(_10103__bF_buf0), .C(_10205_), .Y(_10206_) );
INVX1 INVX1_869 ( .A(_10206_), .Y(_10207_) );
OAI21X1 OAI21X1_2201 ( .A(_10207_), .B(_4431__bF_buf2), .C(_10123__bF_buf1), .Y(_10208_) );
NAND2X1 NAND2X1_638 ( .A(_10167_), .B(_10193_), .Y(_10209_) );
OAI21X1 OAI21X1_2202 ( .A(_10196_), .B(_10190_), .C(_10186_), .Y(_10210_) );
OAI21X1 OAI21X1_2203 ( .A(decoded_imm_uj_5_), .B(_10192_), .C(_10210_), .Y(_10211_) );
OAI21X1 OAI21X1_2204 ( .A(_10188_), .B(_10209_), .C(_10211_), .Y(_10212_) );
INVX1 INVX1_870 ( .A(decoded_imm_uj_6_), .Y(_10213_) );
XNOR2X1 XNOR2X1_19 ( .A(_10206_), .B(_10213_), .Y(_10214_) );
OAI21X1 OAI21X1_2205 ( .A(_10212_), .B(_10214_), .C(instr_jal_bF_buf0), .Y(_10215_) );
AOI21X1 AOI21X1_722 ( .A(_10212_), .B(_10214_), .C(_10215_), .Y(_10216_) );
OR2X2 OR2X2_23 ( .A(_10198_), .B(_10207_), .Y(_10217_) );
OAI21X1 OAI21X1_2206 ( .A(_10180_), .B(_10196_), .C(_10207_), .Y(_10218_) );
NAND2X1 NAND2X1_639 ( .A(_10218_), .B(_10217_), .Y(_10219_) );
OAI21X1 OAI21X1_2207 ( .A(_10219_), .B(instr_jal_bF_buf6), .C(decoder_trigger_bF_buf3), .Y(_10220_) );
OAI21X1 OAI21X1_2208 ( .A(_10216_), .B(_10220_), .C(_10208_), .Y(_10221_) );
AOI21X1 AOI21X1_723 ( .A(_10204_), .B(_10221_), .C(_4426__bF_buf6), .Y(_80__6_) );
NAND2X1 NAND2X1_640 ( .A(reg_next_pc_7_), .B(_4431__bF_buf1), .Y(_10222_) );
NAND2X1 NAND2X1_641 ( .A(_10214_), .B(_10212_), .Y(_10223_) );
OAI21X1 OAI21X1_2209 ( .A(_10213_), .B(_10207_), .C(_10223_), .Y(_10224_) );
INVX1 INVX1_871 ( .A(decoded_imm_uj_7_), .Y(_10225_) );
OAI21X1 OAI21X1_2210 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_7_), .Y(_10226_) );
OAI21X1 OAI21X1_2211 ( .A(_4675_), .B(_10103__bF_buf6), .C(_10226_), .Y(_10227_) );
XNOR2X1 XNOR2X1_20 ( .A(_10227_), .B(_10225_), .Y(_10228_) );
OAI21X1 OAI21X1_2212 ( .A(_10224_), .B(_10228_), .C(instr_jal_bF_buf5), .Y(_10229_) );
AOI21X1 AOI21X1_724 ( .A(_10224_), .B(_10228_), .C(_10229_), .Y(_10230_) );
INVX1 INVX1_872 ( .A(_10227_), .Y(_10231_) );
NOR2X1 NOR2X1_911 ( .A(_10207_), .B(_10231_), .Y(_10232_) );
NAND3X1 NAND3X1_59 ( .A(_10179_), .B(_10197_), .C(_10232_), .Y(_10233_) );
OAI21X1 OAI21X1_2213 ( .A(_10198_), .B(_10207_), .C(_10231_), .Y(_10234_) );
NAND2X1 NAND2X1_642 ( .A(_10233_), .B(_10234_), .Y(_10235_) );
OAI21X1 OAI21X1_2214 ( .A(_10235_), .B(instr_jal_bF_buf4), .C(decoder_trigger_bF_buf2), .Y(_10236_) );
OAI21X1 OAI21X1_2215 ( .A(_10231_), .B(_4431__bF_buf0), .C(_10123__bF_buf0), .Y(_10237_) );
OAI21X1 OAI21X1_2216 ( .A(_10230_), .B(_10236_), .C(_10237_), .Y(_10238_) );
AOI21X1 AOI21X1_725 ( .A(_10222_), .B(_10238_), .C(_4426__bF_buf5), .Y(_80__7_) );
NAND2X1 NAND2X1_643 ( .A(reg_next_pc_8_), .B(_4431__bF_buf7), .Y(_10239_) );
OAI21X1 OAI21X1_2217 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_8_), .Y(_10240_) );
OAI21X1 OAI21X1_2218 ( .A(_4683_), .B(_10103__bF_buf5), .C(_10240_), .Y(_10241_) );
INVX1 INVX1_873 ( .A(_10241_), .Y(_10242_) );
NOR2X1 NOR2X1_912 ( .A(_4431__bF_buf6), .B(_10242_), .Y(_10243_) );
XNOR2X1 XNOR2X1_21 ( .A(_10192_), .B(decoded_imm_uj_5_), .Y(_10244_) );
NOR2X1 NOR2X1_913 ( .A(_10187_), .B(_10244_), .Y(_10245_) );
NAND2X1 NAND2X1_644 ( .A(decoded_imm_uj_6_), .B(_10207_), .Y(_10246_) );
NAND2X1 NAND2X1_645 ( .A(_10213_), .B(_10206_), .Y(_10247_) );
XNOR2X1 XNOR2X1_22 ( .A(_10227_), .B(decoded_imm_uj_7_), .Y(_10248_) );
AOI21X1 AOI21X1_726 ( .A(_10246_), .B(_10247_), .C(_10248_), .Y(_10249_) );
NAND2X1 NAND2X1_646 ( .A(_10249_), .B(_10245_), .Y(_10250_) );
AOI21X1 AOI21X1_727 ( .A(_10170_), .B(_10175_), .C(_10250_), .Y(_10251_) );
NOR2X1 NOR2X1_914 ( .A(_10213_), .B(_10207_), .Y(_10252_) );
NOR2X1 NOR2X1_915 ( .A(_10225_), .B(_10231_), .Y(_10253_) );
AOI21X1 AOI21X1_728 ( .A(_10252_), .B(_10228_), .C(_10253_), .Y(_10254_) );
NAND2X1 NAND2X1_647 ( .A(_10214_), .B(_10228_), .Y(_10255_) );
OAI21X1 OAI21X1_2219 ( .A(_10211_), .B(_10255_), .C(_10254_), .Y(_10256_) );
NOR2X1 NOR2X1_916 ( .A(_10256_), .B(_10251_), .Y(_10257_) );
XNOR2X1 XNOR2X1_23 ( .A(_10241_), .B(decoded_imm_uj_8_), .Y(_10258_) );
OAI21X1 OAI21X1_2220 ( .A(_10257_), .B(_10258_), .C(instr_jal_bF_buf3), .Y(_10259_) );
AOI21X1 AOI21X1_729 ( .A(_10257_), .B(_10258_), .C(_10259_), .Y(_10260_) );
NOR2X1 NOR2X1_917 ( .A(_10242_), .B(_10233_), .Y(_10261_) );
INVX1 INVX1_874 ( .A(_10233_), .Y(_10262_) );
OAI21X1 OAI21X1_2221 ( .A(_10262_), .B(_10241_), .C(_4499__bF_buf0), .Y(_10263_) );
OAI21X1 OAI21X1_2222 ( .A(_10263_), .B(_10261_), .C(decoder_trigger_bF_buf1), .Y(_10264_) );
OAI22X1 OAI22X1_223 ( .A(_10099__bF_buf0), .B(_10243_), .C(_10260_), .D(_10264_), .Y(_10265_) );
AOI21X1 AOI21X1_730 ( .A(_10239_), .B(_10265_), .C(_4426__bF_buf4), .Y(_80__8_) );
NAND2X1 NAND2X1_648 ( .A(reg_next_pc_9_), .B(_4431__bF_buf5), .Y(_10266_) );
NAND2X1 NAND2X1_649 ( .A(decoded_imm_uj_8_), .B(_10241_), .Y(_10267_) );
OAI21X1 OAI21X1_2223 ( .A(_10257_), .B(_10258_), .C(_10267_), .Y(_10268_) );
INVX1 INVX1_875 ( .A(decoded_imm_uj_9_), .Y(_10269_) );
MUX2X1 MUX2X1_208 ( .A(alu_out_q_9_), .B(reg_out_9_), .S(latched_stalu_bF_buf3), .Y(_10270_) );
OAI21X1 OAI21X1_2224 ( .A(_10109__bF_buf1), .B(_4639__bF_buf3), .C(reg_next_pc_9_), .Y(_10271_) );
OAI21X1 OAI21X1_2225 ( .A(_10270_), .B(_10103__bF_buf4), .C(_10271_), .Y(_10272_) );
XNOR2X1 XNOR2X1_24 ( .A(_10272_), .B(_10269_), .Y(_10273_) );
OAI21X1 OAI21X1_2226 ( .A(_10268_), .B(_10273_), .C(instr_jal_bF_buf2), .Y(_10274_) );
AOI21X1 AOI21X1_731 ( .A(_10268_), .B(_10273_), .C(_10274_), .Y(_10275_) );
NAND2X1 NAND2X1_650 ( .A(_10241_), .B(_10272_), .Y(_10276_) );
NOR2X1 NOR2X1_918 ( .A(_10276_), .B(_10233_), .Y(_10277_) );
OAI21X1 OAI21X1_2227 ( .A(_10261_), .B(_10272_), .C(_4499__bF_buf5), .Y(_10278_) );
OAI21X1 OAI21X1_2228 ( .A(_10278_), .B(_10277_), .C(decoder_trigger_bF_buf0), .Y(_10279_) );
MUX2X1 MUX2X1_209 ( .A(_4695_), .B(reg_next_pc_9_), .S(_10118__bF_buf0), .Y(_10280_) );
OAI21X1 OAI21X1_2229 ( .A(_10280_), .B(_4431__bF_buf4), .C(_10123__bF_buf4), .Y(_10281_) );
OAI21X1 OAI21X1_2230 ( .A(_10275_), .B(_10279_), .C(_10281_), .Y(_10282_) );
AOI21X1 AOI21X1_732 ( .A(_10266_), .B(_10282_), .C(_4426__bF_buf3), .Y(_80__9_) );
NAND2X1 NAND2X1_651 ( .A(reg_next_pc_10_), .B(_4431__bF_buf3), .Y(_10283_) );
OAI21X1 OAI21X1_2231 ( .A(_10109__bF_buf0), .B(_4639__bF_buf2), .C(reg_next_pc_10_), .Y(_10284_) );
OAI21X1 OAI21X1_2232 ( .A(_4698_), .B(_10103__bF_buf3), .C(_10284_), .Y(_10285_) );
INVX1 INVX1_876 ( .A(_10285_), .Y(_10286_) );
OAI21X1 OAI21X1_2233 ( .A(_10286_), .B(_4431__bF_buf2), .C(_10123__bF_buf3), .Y(_10287_) );
INVX1 INVX1_877 ( .A(decoded_imm_uj_10_), .Y(_10288_) );
XNOR2X1 XNOR2X1_25 ( .A(_10285_), .B(_10288_), .Y(_10289_) );
NAND2X1 NAND2X1_652 ( .A(decoded_imm_uj_5_), .B(_10192_), .Y(_10290_) );
OAI21X1 OAI21X1_2234 ( .A(_10244_), .B(_10186_), .C(_10290_), .Y(_10291_) );
OAI21X1 OAI21X1_2235 ( .A(decoded_imm_uj_7_), .B(_10227_), .C(_10252_), .Y(_10292_) );
OAI21X1 OAI21X1_2236 ( .A(_10225_), .B(_10231_), .C(_10292_), .Y(_10293_) );
AOI21X1 AOI21X1_733 ( .A(_10249_), .B(_10291_), .C(_10293_), .Y(_10294_) );
OAI21X1 OAI21X1_2237 ( .A(_10188_), .B(_10250_), .C(_10294_), .Y(_10295_) );
XNOR2X1 XNOR2X1_26 ( .A(_10272_), .B(decoded_imm_uj_9_), .Y(_10296_) );
NOR2X1 NOR2X1_919 ( .A(_10258_), .B(_10296_), .Y(_10297_) );
OAI21X1 OAI21X1_2238 ( .A(_10269_), .B(_10280_), .C(_10267_), .Y(_10298_) );
OAI21X1 OAI21X1_2239 ( .A(decoded_imm_uj_9_), .B(_10272_), .C(_10298_), .Y(_10299_) );
INVX1 INVX1_878 ( .A(_10299_), .Y(_10300_) );
AOI21X1 AOI21X1_734 ( .A(_10297_), .B(_10295_), .C(_10300_), .Y(_10301_) );
INVX1 INVX1_879 ( .A(_10301_), .Y(_10302_) );
OAI21X1 OAI21X1_2240 ( .A(_10302_), .B(_10289_), .C(instr_jal_bF_buf1), .Y(_10303_) );
AOI21X1 AOI21X1_735 ( .A(_10289_), .B(_10302_), .C(_10303_), .Y(_10304_) );
NAND2X1 NAND2X1_653 ( .A(_10285_), .B(_10277_), .Y(_10305_) );
OAI21X1 OAI21X1_2241 ( .A(_10233_), .B(_10276_), .C(_10286_), .Y(_10306_) );
NAND2X1 NAND2X1_654 ( .A(_10306_), .B(_10305_), .Y(_10307_) );
OAI21X1 OAI21X1_2242 ( .A(_10307_), .B(instr_jal_bF_buf0), .C(decoder_trigger_bF_buf3), .Y(_10308_) );
OAI21X1 OAI21X1_2243 ( .A(_10304_), .B(_10308_), .C(_10287_), .Y(_10309_) );
AOI21X1 AOI21X1_736 ( .A(_10283_), .B(_10309_), .C(_4426__bF_buf2), .Y(_80__10_) );
NAND2X1 NAND2X1_655 ( .A(reg_next_pc_11_), .B(_4431__bF_buf1), .Y(_10310_) );
NAND2X1 NAND2X1_656 ( .A(_10289_), .B(_10302_), .Y(_10311_) );
OAI21X1 OAI21X1_2244 ( .A(_10288_), .B(_10286_), .C(_10311_), .Y(_10312_) );
INVX1 INVX1_880 ( .A(decoded_imm_uj_11_), .Y(_10313_) );
OAI21X1 OAI21X1_2245 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_11_), .Y(_10314_) );
OAI21X1 OAI21X1_2246 ( .A(_4705_), .B(_10103__bF_buf2), .C(_10314_), .Y(_10315_) );
XNOR2X1 XNOR2X1_27 ( .A(_10315_), .B(_10313_), .Y(_10316_) );
AOI21X1 AOI21X1_737 ( .A(_10316_), .B(_10312_), .C(_4499__bF_buf4), .Y(_10317_) );
OAI21X1 OAI21X1_2247 ( .A(_10312_), .B(_10316_), .C(_10317_), .Y(_10318_) );
INVX1 INVX1_881 ( .A(_10315_), .Y(_10319_) );
NAND2X1 NAND2X1_657 ( .A(_10319_), .B(_10305_), .Y(_10320_) );
NAND2X1 NAND2X1_658 ( .A(_10285_), .B(_10315_), .Y(_10321_) );
NOR2X1 NOR2X1_920 ( .A(_10276_), .B(_10321_), .Y(_10322_) );
INVX1 INVX1_882 ( .A(_10322_), .Y(_10323_) );
OR2X2 OR2X2_24 ( .A(_10233_), .B(_10323_), .Y(_10324_) );
AOI21X1 AOI21X1_738 ( .A(_10324_), .B(_10320_), .C(_4605__bF_buf1), .Y(_10325_) );
OAI21X1 OAI21X1_2248 ( .A(_10107_), .B(_10325_), .C(_10318_), .Y(_10326_) );
NOR2X1 NOR2X1_921 ( .A(_4431__bF_buf0), .B(_10319_), .Y(_10327_) );
OAI21X1 OAI21X1_2249 ( .A(_10099__bF_buf3), .B(_10327_), .C(_10326_), .Y(_10328_) );
AOI21X1 AOI21X1_739 ( .A(_10310_), .B(_10328_), .C(_4426__bF_buf1), .Y(_80__11_) );
NAND2X1 NAND2X1_659 ( .A(reg_next_pc_12_), .B(_4431__bF_buf7), .Y(_10329_) );
OAI21X1 OAI21X1_2250 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_12_), .Y(_10330_) );
OAI21X1 OAI21X1_2251 ( .A(_4716_), .B(_10103__bF_buf1), .C(_10330_), .Y(_10331_) );
NAND2X1 NAND2X1_660 ( .A(cpu_state_1_bF_buf3_), .B(_10331_), .Y(_10332_) );
OAI21X1 OAI21X1_2252 ( .A(_4431__bF_buf6), .B(_4605__bF_buf0), .C(_10332_), .Y(_10333_) );
NOR2X1 NOR2X1_922 ( .A(_10288_), .B(_10286_), .Y(_10334_) );
NOR2X1 NOR2X1_923 ( .A(_10313_), .B(_10319_), .Y(_10335_) );
AOI21X1 AOI21X1_740 ( .A(_10334_), .B(_10316_), .C(_10335_), .Y(_10336_) );
NAND2X1 NAND2X1_661 ( .A(_10289_), .B(_10316_), .Y(_10337_) );
OAI21X1 OAI21X1_2253 ( .A(_10299_), .B(_10337_), .C(_10336_), .Y(_10338_) );
INVX1 INVX1_883 ( .A(decoded_imm_uj_8_), .Y(_10339_) );
XNOR2X1 XNOR2X1_28 ( .A(_10241_), .B(_10339_), .Y(_10340_) );
NAND2X1 NAND2X1_662 ( .A(_10340_), .B(_10273_), .Y(_10341_) );
NOR2X1 NOR2X1_924 ( .A(_10341_), .B(_10337_), .Y(_10342_) );
AOI21X1 AOI21X1_741 ( .A(_10342_), .B(_10295_), .C(_10338_), .Y(_10343_) );
XNOR2X1 XNOR2X1_29 ( .A(_10331_), .B(decoded_imm_uj_12_), .Y(_10344_) );
NOR2X1 NOR2X1_925 ( .A(_10344_), .B(_10343_), .Y(_10345_) );
INVX1 INVX1_884 ( .A(_10343_), .Y(_10346_) );
INVX1 INVX1_885 ( .A(decoded_imm_uj_12_), .Y(_10347_) );
XNOR2X1 XNOR2X1_30 ( .A(_10331_), .B(_10347_), .Y(_10348_) );
OAI21X1 OAI21X1_2254 ( .A(_10346_), .B(_10348_), .C(instr_jal_bF_buf6), .Y(_10349_) );
NOR2X1 NOR2X1_926 ( .A(_10345_), .B(_10349_), .Y(_10350_) );
INVX1 INVX1_886 ( .A(_10324_), .Y(_10351_) );
NAND2X1 NAND2X1_663 ( .A(_10331_), .B(_10351_), .Y(_10352_) );
INVX1 INVX1_887 ( .A(_10331_), .Y(_10353_) );
OAI21X1 OAI21X1_2255 ( .A(_10233_), .B(_10323_), .C(_10353_), .Y(_10354_) );
NAND2X1 NAND2X1_664 ( .A(_10354_), .B(_10352_), .Y(_10355_) );
OAI21X1 OAI21X1_2256 ( .A(_10355_), .B(instr_jal_bF_buf5), .C(decoder_trigger_bF_buf2), .Y(_10356_) );
OAI21X1 OAI21X1_2257 ( .A(_10350_), .B(_10356_), .C(_10333_), .Y(_10357_) );
AOI21X1 AOI21X1_742 ( .A(_10329_), .B(_10357_), .C(_4426__bF_buf0), .Y(_80__12_) );
NAND2X1 NAND2X1_665 ( .A(reg_next_pc_13_), .B(_4431__bF_buf5), .Y(_10358_) );
AOI21X1 AOI21X1_743 ( .A(decoded_imm_uj_12_), .B(_10331_), .C(_10345_), .Y(_10359_) );
INVX1 INVX1_888 ( .A(decoded_imm_uj_13_), .Y(_10360_) );
MUX2X1 MUX2X1_210 ( .A(_4726_), .B(reg_next_pc_13_), .S(_10118__bF_buf4), .Y(_10361_) );
NAND2X1 NAND2X1_666 ( .A(_10360_), .B(_10361_), .Y(_10362_) );
MUX2X1 MUX2X1_211 ( .A(alu_out_q_13_), .B(reg_out_13_), .S(latched_stalu_bF_buf2), .Y(_10363_) );
OAI21X1 OAI21X1_2258 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_13_), .Y(_10364_) );
OAI21X1 OAI21X1_2259 ( .A(_10363_), .B(_10103__bF_buf0), .C(_10364_), .Y(_10365_) );
NAND2X1 NAND2X1_667 ( .A(decoded_imm_uj_13_), .B(_10365_), .Y(_10366_) );
NAND2X1 NAND2X1_668 ( .A(_10366_), .B(_10362_), .Y(_10367_) );
AND2X2 AND2X2_163 ( .A(_10359_), .B(_10367_), .Y(_10368_) );
OAI21X1 OAI21X1_2260 ( .A(_10359_), .B(_10367_), .C(instr_jal_bF_buf4), .Y(_10369_) );
OAI21X1 OAI21X1_2261 ( .A(_10324_), .B(_10353_), .C(_10361_), .Y(_10370_) );
NAND2X1 NAND2X1_669 ( .A(_10331_), .B(_10365_), .Y(_10371_) );
OR2X2 OR2X2_25 ( .A(_10324_), .B(_10371_), .Y(_10372_) );
AOI21X1 AOI21X1_744 ( .A(_10370_), .B(_10372_), .C(_4605__bF_buf5), .Y(_10373_) );
OAI22X1 OAI22X1_224 ( .A(_10107_), .B(_10373_), .C(_10368_), .D(_10369_), .Y(_10374_) );
NOR2X1 NOR2X1_927 ( .A(_4431__bF_buf4), .B(_10361_), .Y(_10375_) );
OAI21X1 OAI21X1_2262 ( .A(_10099__bF_buf2), .B(_10375_), .C(_10374_), .Y(_10376_) );
AOI21X1 AOI21X1_745 ( .A(_10358_), .B(_10376_), .C(_4426__bF_buf11), .Y(_80__13_) );
NAND2X1 NAND2X1_670 ( .A(reg_next_pc_14_), .B(_4431__bF_buf3), .Y(_10377_) );
OAI21X1 OAI21X1_2263 ( .A(_10109__bF_buf1), .B(_4639__bF_buf3), .C(reg_next_pc_14_), .Y(_10378_) );
OAI21X1 OAI21X1_2264 ( .A(_4733_), .B(_10103__bF_buf6), .C(_10378_), .Y(_10379_) );
INVX1 INVX1_889 ( .A(_10379_), .Y(_10380_) );
OAI21X1 OAI21X1_2265 ( .A(_10380_), .B(_4431__bF_buf2), .C(_10123__bF_buf2), .Y(_10381_) );
INVX1 INVX1_890 ( .A(decoded_imm_uj_14_), .Y(_10382_) );
XNOR2X1 XNOR2X1_31 ( .A(_10379_), .B(_10382_), .Y(_10383_) );
NAND2X1 NAND2X1_671 ( .A(decoded_imm_uj_12_), .B(_10331_), .Y(_10384_) );
OAI21X1 OAI21X1_2266 ( .A(_10360_), .B(_10361_), .C(_10384_), .Y(_10385_) );
OAI21X1 OAI21X1_2267 ( .A(decoded_imm_uj_13_), .B(_10365_), .C(_10385_), .Y(_10386_) );
NAND3X1 NAND3X1_60 ( .A(_10362_), .B(_10366_), .C(_10348_), .Y(_10387_) );
OAI21X1 OAI21X1_2268 ( .A(_10343_), .B(_10387_), .C(_10386_), .Y(_10388_) );
NAND2X1 NAND2X1_672 ( .A(_10383_), .B(_10388_), .Y(_10389_) );
INVX1 INVX1_891 ( .A(_10389_), .Y(_10390_) );
XNOR2X1 XNOR2X1_32 ( .A(_10372_), .B(_10380_), .Y(_10391_) );
OAI21X1 OAI21X1_2269 ( .A(_10388_), .B(_10383_), .C(instr_jal_bF_buf3), .Y(_10392_) );
OAI22X1 OAI22X1_225 ( .A(instr_jal_bF_buf2), .B(_10391_), .C(_10390_), .D(_10392_), .Y(_10393_) );
OAI21X1 OAI21X1_2270 ( .A(_10393_), .B(_4605__bF_buf4), .C(_10381_), .Y(_10394_) );
AOI21X1 AOI21X1_746 ( .A(_10377_), .B(_10394_), .C(_4426__bF_buf10), .Y(_80__14_) );
NAND2X1 NAND2X1_673 ( .A(reg_next_pc_15_), .B(_4431__bF_buf1), .Y(_10395_) );
OAI21X1 OAI21X1_2271 ( .A(_10382_), .B(_10380_), .C(_10389_), .Y(_10396_) );
INVX1 INVX1_892 ( .A(decoded_imm_uj_15_), .Y(_10397_) );
OAI21X1 OAI21X1_2272 ( .A(_10109__bF_buf0), .B(_4639__bF_buf2), .C(reg_next_pc_15_), .Y(_10398_) );
OAI21X1 OAI21X1_2273 ( .A(_4742_), .B(_10103__bF_buf5), .C(_10398_), .Y(_10399_) );
XNOR2X1 XNOR2X1_33 ( .A(_10399_), .B(_10397_), .Y(_10400_) );
OAI21X1 OAI21X1_2274 ( .A(_10396_), .B(_10400_), .C(instr_jal_bF_buf1), .Y(_10401_) );
AOI21X1 AOI21X1_747 ( .A(_10396_), .B(_10400_), .C(_10401_), .Y(_10402_) );
INVX1 INVX1_893 ( .A(_10399_), .Y(_10403_) );
OAI21X1 OAI21X1_2275 ( .A(_10372_), .B(_10380_), .C(_10403_), .Y(_10404_) );
INVX1 INVX1_894 ( .A(_10378_), .Y(_10405_) );
NOR2X1 NOR2X1_928 ( .A(_10103__bF_buf4), .B(_4733_), .Y(_10406_) );
OAI21X1 OAI21X1_2276 ( .A(_10406_), .B(_10405_), .C(_10399_), .Y(_10407_) );
OR2X2 OR2X2_26 ( .A(_10407_), .B(_10361_), .Y(_10408_) );
OAI21X1 OAI21X1_2277 ( .A(_10352_), .B(_10408_), .C(_10404_), .Y(_10409_) );
OAI21X1 OAI21X1_2278 ( .A(_10409_), .B(instr_jal_bF_buf0), .C(decoder_trigger_bF_buf1), .Y(_10410_) );
OAI21X1 OAI21X1_2279 ( .A(_10403_), .B(_4431__bF_buf0), .C(_10123__bF_buf1), .Y(_10411_) );
OAI21X1 OAI21X1_2280 ( .A(_10402_), .B(_10410_), .C(_10411_), .Y(_10412_) );
AOI21X1 AOI21X1_748 ( .A(_10395_), .B(_10412_), .C(_4426__bF_buf9), .Y(_80__15_) );
NAND2X1 NAND2X1_674 ( .A(reg_next_pc_16_), .B(_4431__bF_buf7), .Y(_10413_) );
MUX2X1 MUX2X1_212 ( .A(_4751_), .B(reg_next_pc_16_), .S(_10118__bF_buf3), .Y(_10414_) );
OAI21X1 OAI21X1_2281 ( .A(_10414_), .B(_4431__bF_buf6), .C(_10123__bF_buf0), .Y(_10415_) );
NAND3X1 NAND3X1_61 ( .A(_10289_), .B(_10316_), .C(_10297_), .Y(_10416_) );
NOR2X1 NOR2X1_929 ( .A(_10344_), .B(_10367_), .Y(_10417_) );
AND2X2 AND2X2_164 ( .A(_10383_), .B(_10400_), .Y(_10418_) );
NAND2X1 NAND2X1_675 ( .A(_10417_), .B(_10418_), .Y(_10419_) );
NOR2X1 NOR2X1_930 ( .A(_10419_), .B(_10416_), .Y(_10420_) );
OAI21X1 OAI21X1_2282 ( .A(_10251_), .B(_10256_), .C(_10420_), .Y(_10421_) );
NAND2X1 NAND2X1_676 ( .A(_10383_), .B(_10400_), .Y(_10422_) );
NOR2X1 NOR2X1_931 ( .A(_10422_), .B(_10387_), .Y(_10423_) );
NOR2X1 NOR2X1_932 ( .A(_10382_), .B(_10380_), .Y(_10424_) );
NOR2X1 NOR2X1_933 ( .A(_10397_), .B(_10403_), .Y(_10425_) );
AOI21X1 AOI21X1_749 ( .A(_10424_), .B(_10400_), .C(_10425_), .Y(_10426_) );
OAI21X1 OAI21X1_2283 ( .A(_10386_), .B(_10422_), .C(_10426_), .Y(_10427_) );
AOI21X1 AOI21X1_750 ( .A(_10423_), .B(_10338_), .C(_10427_), .Y(_10428_) );
OAI21X1 OAI21X1_2284 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_16_), .Y(_10429_) );
NAND2X1 NAND2X1_677 ( .A(_10118__bF_buf2), .B(_4751_), .Y(_10430_) );
NAND2X1 NAND2X1_678 ( .A(_10429_), .B(_10430_), .Y(_10431_) );
NAND2X1 NAND2X1_679 ( .A(decoded_imm_uj_16_), .B(_10431_), .Y(_10432_) );
INVX1 INVX1_895 ( .A(decoded_imm_uj_16_), .Y(_10433_) );
NAND2X1 NAND2X1_680 ( .A(_10433_), .B(_10414_), .Y(_10434_) );
AND2X2 AND2X2_165 ( .A(_10432_), .B(_10434_), .Y(_10435_) );
INVX1 INVX1_896 ( .A(_10435_), .Y(_10436_) );
AOI21X1 AOI21X1_751 ( .A(_10428_), .B(_10421_), .C(_10436_), .Y(_10437_) );
NAND2X1 NAND2X1_681 ( .A(_10342_), .B(_10423_), .Y(_10438_) );
OAI21X1 OAI21X1_2285 ( .A(_10257_), .B(_10438_), .C(_10428_), .Y(_10439_) );
OAI21X1 OAI21X1_2286 ( .A(_10439_), .B(_10435_), .C(instr_jal_bF_buf6), .Y(_10440_) );
NOR2X1 NOR2X1_934 ( .A(_10437_), .B(_10440_), .Y(_10441_) );
NOR3X1 NOR3X1_2 ( .A(_10353_), .B(_10408_), .C(_10324_), .Y(_10442_) );
AND2X2 AND2X2_166 ( .A(_10442_), .B(_10431_), .Y(_10443_) );
OAI21X1 OAI21X1_2287 ( .A(_10442_), .B(_10431_), .C(_4499__bF_buf3), .Y(_10444_) );
OAI21X1 OAI21X1_2288 ( .A(_10443_), .B(_10444_), .C(decoder_trigger_bF_buf0), .Y(_10445_) );
OAI21X1 OAI21X1_2289 ( .A(_10441_), .B(_10445_), .C(_10415_), .Y(_10446_) );
AOI21X1 AOI21X1_752 ( .A(_10413_), .B(_10446_), .C(_4426__bF_buf8), .Y(_80__16_) );
NAND2X1 NAND2X1_682 ( .A(reg_next_pc_17_), .B(_4431__bF_buf5), .Y(_10447_) );
INVX1 INVX1_897 ( .A(_10437_), .Y(_10448_) );
OAI21X1 OAI21X1_2290 ( .A(_10433_), .B(_10414_), .C(_10448_), .Y(_10449_) );
OAI21X1 OAI21X1_2291 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_17_), .Y(_10450_) );
NAND2X1 NAND2X1_683 ( .A(_10118__bF_buf1), .B(_4759_), .Y(_10451_) );
NAND2X1 NAND2X1_684 ( .A(_10450_), .B(_10451_), .Y(_10452_) );
NAND2X1 NAND2X1_685 ( .A(decoded_imm_uj_17_), .B(_10452_), .Y(_10453_) );
INVX1 INVX1_898 ( .A(decoded_imm_uj_17_), .Y(_10454_) );
MUX2X1 MUX2X1_213 ( .A(_4759_), .B(reg_next_pc_17_), .S(_10118__bF_buf0), .Y(_10455_) );
NAND2X1 NAND2X1_686 ( .A(_10454_), .B(_10455_), .Y(_10456_) );
AND2X2 AND2X2_167 ( .A(_10453_), .B(_10456_), .Y(_10457_) );
OAI21X1 OAI21X1_2292 ( .A(_10449_), .B(_10457_), .C(instr_jal_bF_buf5), .Y(_10458_) );
AOI21X1 AOI21X1_753 ( .A(_10449_), .B(_10457_), .C(_10458_), .Y(_10459_) );
NOR2X1 NOR2X1_935 ( .A(_10452_), .B(_10443_), .Y(_10460_) );
NOR2X1 NOR2X1_936 ( .A(_10414_), .B(_10455_), .Y(_10461_) );
NAND2X1 NAND2X1_687 ( .A(_10461_), .B(_10442_), .Y(_10462_) );
NAND2X1 NAND2X1_688 ( .A(_4499__bF_buf2), .B(_10462_), .Y(_10463_) );
OAI21X1 OAI21X1_2293 ( .A(_10460_), .B(_10463_), .C(decoder_trigger_bF_buf3), .Y(_10464_) );
NOR2X1 NOR2X1_937 ( .A(_4431__bF_buf4), .B(_10455_), .Y(_10465_) );
OAI22X1 OAI22X1_226 ( .A(_10099__bF_buf1), .B(_10465_), .C(_10459_), .D(_10464_), .Y(_10466_) );
AOI21X1 AOI21X1_754 ( .A(_10447_), .B(_10466_), .C(_4426__bF_buf7), .Y(_80__17_) );
NAND2X1 NAND2X1_689 ( .A(reg_next_pc_18_), .B(_4431__bF_buf3), .Y(_10467_) );
MUX2X1 MUX2X1_214 ( .A(_4767_), .B(reg_next_pc_18_), .S(_10118__bF_buf4), .Y(_10468_) );
OAI21X1 OAI21X1_2294 ( .A(_10468_), .B(_4431__bF_buf2), .C(_10123__bF_buf4), .Y(_10469_) );
INVX1 INVX1_899 ( .A(decoded_imm_uj_18_), .Y(_10470_) );
NOR2X1 NOR2X1_938 ( .A(_10470_), .B(_10468_), .Y(_10471_) );
OAI21X1 OAI21X1_2295 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_18_), .Y(_10472_) );
NAND2X1 NAND2X1_690 ( .A(_10118__bF_buf3), .B(_4767_), .Y(_10473_) );
NAND2X1 NAND2X1_691 ( .A(_10472_), .B(_10473_), .Y(_10474_) );
NOR2X1 NOR2X1_939 ( .A(decoded_imm_uj_18_), .B(_10474_), .Y(_10475_) );
NOR2X1 NOR2X1_940 ( .A(_10471_), .B(_10475_), .Y(_10476_) );
OAI21X1 OAI21X1_2296 ( .A(_10433_), .B(_10414_), .C(_10453_), .Y(_10477_) );
OAI21X1 OAI21X1_2297 ( .A(_10437_), .B(_10477_), .C(_10456_), .Y(_10478_) );
NAND2X1 NAND2X1_692 ( .A(_10476_), .B(_10478_), .Y(_10479_) );
OR2X2 OR2X2_27 ( .A(_10478_), .B(_10476_), .Y(_10480_) );
AOI21X1 AOI21X1_755 ( .A(_10479_), .B(_10480_), .C(_4499__bF_buf1), .Y(_10481_) );
NAND3X1 NAND3X1_62 ( .A(_10461_), .B(_10474_), .C(_10442_), .Y(_10482_) );
NAND2X1 NAND2X1_693 ( .A(_10468_), .B(_10462_), .Y(_10483_) );
NAND2X1 NAND2X1_694 ( .A(_10482_), .B(_10483_), .Y(_10484_) );
OAI21X1 OAI21X1_2298 ( .A(_10484_), .B(instr_jal_bF_buf4), .C(decoder_trigger_bF_buf2), .Y(_10485_) );
OAI21X1 OAI21X1_2299 ( .A(_10481_), .B(_10485_), .C(_10469_), .Y(_10486_) );
AOI21X1 AOI21X1_756 ( .A(_10467_), .B(_10486_), .C(_4426__bF_buf6), .Y(_80__18_) );
INVX1 INVX1_900 ( .A(reg_next_pc_19_), .Y(_10487_) );
INVX1 INVX1_901 ( .A(_10471_), .Y(_10488_) );
OAI21X1 OAI21X1_2300 ( .A(_10478_), .B(_10475_), .C(_10488_), .Y(_10489_) );
INVX1 INVX1_902 ( .A(decoded_imm_uj_19_), .Y(_10490_) );
NOR2X1 NOR2X1_941 ( .A(_10487_), .B(_10118__bF_buf2), .Y(_10491_) );
AOI21X1 AOI21X1_757 ( .A(_10118__bF_buf1), .B(_4787_), .C(_10491_), .Y(_10492_) );
NOR2X1 NOR2X1_942 ( .A(_10490_), .B(_10492_), .Y(_10493_) );
NAND2X1 NAND2X1_695 ( .A(_10118__bF_buf0), .B(_4787_), .Y(_10494_) );
OAI21X1 OAI21X1_2301 ( .A(_10487_), .B(_10118__bF_buf4), .C(_10494_), .Y(_10495_) );
NOR2X1 NOR2X1_943 ( .A(decoded_imm_uj_19_), .B(_10495_), .Y(_10496_) );
NOR2X1 NOR2X1_944 ( .A(_10493_), .B(_10496_), .Y(_10497_) );
OAI21X1 OAI21X1_2302 ( .A(_10489_), .B(_10497_), .C(instr_jal_bF_buf3), .Y(_10498_) );
AOI21X1 AOI21X1_758 ( .A(_10489_), .B(_10497_), .C(_10498_), .Y(_10499_) );
OAI21X1 OAI21X1_2303 ( .A(_10462_), .B(_10468_), .C(_10492_), .Y(_10500_) );
OR2X2 OR2X2_28 ( .A(_10482_), .B(_10492_), .Y(_10501_) );
NAND2X1 NAND2X1_696 ( .A(_10500_), .B(_10501_), .Y(_10502_) );
OAI21X1 OAI21X1_2304 ( .A(_10502_), .B(instr_jal_bF_buf2), .C(decoder_trigger_bF_buf1), .Y(_10503_) );
OAI21X1 OAI21X1_2305 ( .A(_10492_), .B(_4431__bF_buf1), .C(_10123__bF_buf3), .Y(_10504_) );
OAI21X1 OAI21X1_2306 ( .A(_10499_), .B(_10503_), .C(_10504_), .Y(_10505_) );
OAI21X1 OAI21X1_2307 ( .A(cpu_state_1_bF_buf2_), .B(_10487_), .C(_10505_), .Y(_10506_) );
AND2X2 AND2X2_168 ( .A(_10506_), .B(resetn_bF_buf1), .Y(_80__19_) );
NAND2X1 NAND2X1_697 ( .A(reg_next_pc_20_), .B(_4431__bF_buf0), .Y(_10507_) );
MUX2X1 MUX2X1_215 ( .A(_4797_), .B(reg_next_pc_20_), .S(_10118__bF_buf3), .Y(_10508_) );
NOR2X1 NOR2X1_945 ( .A(_4431__bF_buf7), .B(_10508_), .Y(_10509_) );
OAI21X1 OAI21X1_2308 ( .A(decoded_imm_uj_17_), .B(_10452_), .C(_10477_), .Y(_10510_) );
NAND2X1 NAND2X1_698 ( .A(_10476_), .B(_10497_), .Y(_10511_) );
AOI21X1 AOI21X1_759 ( .A(_10471_), .B(_10497_), .C(_10493_), .Y(_10512_) );
OAI21X1 OAI21X1_2309 ( .A(_10510_), .B(_10511_), .C(_10512_), .Y(_10513_) );
NAND2X1 NAND2X1_699 ( .A(_10457_), .B(_10435_), .Y(_10514_) );
NOR2X1 NOR2X1_946 ( .A(_10514_), .B(_10511_), .Y(_10515_) );
AOI21X1 AOI21X1_760 ( .A(_10515_), .B(_10439_), .C(_10513_), .Y(_10516_) );
INVX1 INVX1_903 ( .A(_10508_), .Y(_10517_) );
NAND2X1 NAND2X1_700 ( .A(decoded_imm_uj_20_), .B(_10517_), .Y(_10518_) );
INVX1 INVX1_904 ( .A(decoded_imm_uj_20_), .Y(_10519_) );
NAND2X1 NAND2X1_701 ( .A(_10519_), .B(_10508_), .Y(_10520_) );
AND2X2 AND2X2_169 ( .A(_10518_), .B(_10520_), .Y(_10521_) );
INVX1 INVX1_905 ( .A(_10521_), .Y(_10522_) );
AND2X2 AND2X2_170 ( .A(_10516_), .B(_10522_), .Y(_10523_) );
OAI21X1 OAI21X1_2310 ( .A(_10516_), .B(_10522_), .C(instr_jal_bF_buf1), .Y(_10524_) );
NOR2X1 NOR2X1_947 ( .A(_10371_), .B(_10407_), .Y(_10525_) );
NAND2X1 NAND2X1_702 ( .A(_10322_), .B(_10525_), .Y(_10526_) );
NOR2X1 NOR2X1_948 ( .A(_10233_), .B(_10526_), .Y(_10527_) );
INVX1 INVX1_906 ( .A(_10527_), .Y(_10528_) );
NAND3X1 NAND3X1_63 ( .A(_10474_), .B(_10495_), .C(_10461_), .Y(_10529_) );
NOR2X1 NOR2X1_949 ( .A(_10529_), .B(_10528_), .Y(_10530_) );
XNOR2X1 XNOR2X1_34 ( .A(_10530_), .B(_10508_), .Y(_10531_) );
AOI21X1 AOI21X1_761 ( .A(_4499__bF_buf0), .B(_10531_), .C(_4605__bF_buf3), .Y(_10532_) );
OAI21X1 OAI21X1_2311 ( .A(_10523_), .B(_10524_), .C(_10532_), .Y(_10533_) );
OAI21X1 OAI21X1_2312 ( .A(_10099__bF_buf0), .B(_10509_), .C(_10533_), .Y(_10534_) );
AOI21X1 AOI21X1_762 ( .A(_10507_), .B(_10534_), .C(_4426__bF_buf5), .Y(_80__20_) );
INVX1 INVX1_907 ( .A(reg_next_pc_21_), .Y(_10535_) );
OAI21X1 OAI21X1_2313 ( .A(_10516_), .B(_10522_), .C(_10518_), .Y(_10536_) );
INVX1 INVX1_908 ( .A(decoded_imm_uj_21_), .Y(_10537_) );
NOR2X1 NOR2X1_950 ( .A(_10535_), .B(_10118__bF_buf2), .Y(_10538_) );
AOI21X1 AOI21X1_763 ( .A(_10118__bF_buf1), .B(_4810_), .C(_10538_), .Y(_10539_) );
NOR2X1 NOR2X1_951 ( .A(_10537_), .B(_10539_), .Y(_10540_) );
INVX1 INVX1_909 ( .A(_4810_), .Y(_10541_) );
INVX1 INVX1_910 ( .A(_10538_), .Y(_10542_) );
OAI21X1 OAI21X1_2314 ( .A(_10541_), .B(_10103__bF_buf3), .C(_10542_), .Y(_10543_) );
NOR2X1 NOR2X1_952 ( .A(decoded_imm_uj_21_), .B(_10543_), .Y(_10544_) );
NOR2X1 NOR2X1_953 ( .A(_10540_), .B(_10544_), .Y(_10545_) );
OAI21X1 OAI21X1_2315 ( .A(_10536_), .B(_10545_), .C(instr_jal_bF_buf0), .Y(_10546_) );
AOI21X1 AOI21X1_764 ( .A(_10536_), .B(_10545_), .C(_10546_), .Y(_10547_) );
AOI21X1 AOI21X1_765 ( .A(_10517_), .B(_10530_), .C(_10539_), .Y(_10548_) );
NAND2X1 NAND2X1_703 ( .A(_10517_), .B(_10530_), .Y(_10549_) );
NOR2X1 NOR2X1_954 ( .A(_10543_), .B(_10549_), .Y(_10550_) );
OAI21X1 OAI21X1_2316 ( .A(_10550_), .B(_10548_), .C(_4499__bF_buf5), .Y(_10551_) );
NAND2X1 NAND2X1_704 ( .A(decoder_trigger_bF_buf0), .B(_10551_), .Y(_10552_) );
OAI21X1 OAI21X1_2317 ( .A(_10539_), .B(_4431__bF_buf6), .C(_10123__bF_buf2), .Y(_10553_) );
OAI21X1 OAI21X1_2318 ( .A(_10547_), .B(_10552_), .C(_10553_), .Y(_10554_) );
OAI21X1 OAI21X1_2319 ( .A(cpu_state_1_bF_buf1_), .B(_10535_), .C(_10554_), .Y(_10555_) );
AND2X2 AND2X2_171 ( .A(_10555_), .B(resetn_bF_buf0), .Y(_80__21_) );
NAND2X1 NAND2X1_705 ( .A(reg_next_pc_22_), .B(_4431__bF_buf5), .Y(_10556_) );
MUX2X1 MUX2X1_216 ( .A(_4820_), .B(reg_next_pc_22_), .S(_10118__bF_buf0), .Y(_10557_) );
OAI21X1 OAI21X1_2320 ( .A(_10557_), .B(_4431__bF_buf4), .C(_10123__bF_buf1), .Y(_10558_) );
INVX1 INVX1_911 ( .A(decoded_imm_uj_22_), .Y(_10559_) );
NOR2X1 NOR2X1_955 ( .A(_10559_), .B(_10557_), .Y(_10560_) );
INVX1 INVX1_912 ( .A(_10557_), .Y(_10561_) );
NOR2X1 NOR2X1_956 ( .A(decoded_imm_uj_22_), .B(_10561_), .Y(_10562_) );
NOR2X1 NOR2X1_957 ( .A(_10560_), .B(_10562_), .Y(_10563_) );
NOR2X1 NOR2X1_958 ( .A(_10518_), .B(_10544_), .Y(_10564_) );
NOR2X1 NOR2X1_959 ( .A(_10540_), .B(_10564_), .Y(_10565_) );
NAND2X1 NAND2X1_706 ( .A(_10521_), .B(_10545_), .Y(_10566_) );
OAI21X1 OAI21X1_2321 ( .A(_10516_), .B(_10566_), .C(_10565_), .Y(_10567_) );
AND2X2 AND2X2_172 ( .A(_10567_), .B(_10563_), .Y(_10568_) );
OAI21X1 OAI21X1_2322 ( .A(_10567_), .B(_10563_), .C(instr_jal_bF_buf6), .Y(_10569_) );
NOR2X1 NOR2X1_960 ( .A(_10508_), .B(_10539_), .Y(_10570_) );
AND2X2 AND2X2_173 ( .A(_10530_), .B(_10570_), .Y(_10571_) );
NOR2X1 NOR2X1_961 ( .A(_10557_), .B(_10571_), .Y(_10572_) );
AND2X2 AND2X2_174 ( .A(_10571_), .B(_10557_), .Y(_10573_) );
OAI21X1 OAI21X1_2323 ( .A(_10573_), .B(_10572_), .C(_4499__bF_buf4), .Y(_10574_) );
OAI21X1 OAI21X1_2324 ( .A(_10568_), .B(_10569_), .C(_10574_), .Y(_10575_) );
OAI21X1 OAI21X1_2325 ( .A(_10575_), .B(_4605__bF_buf2), .C(_10558_), .Y(_10576_) );
AOI21X1 AOI21X1_766 ( .A(_10556_), .B(_10576_), .C(_4426__bF_buf4), .Y(_80__22_) );
NAND2X1 NAND2X1_707 ( .A(reg_next_pc_23_), .B(_4431__bF_buf3), .Y(_10577_) );
AOI21X1 AOI21X1_767 ( .A(_10563_), .B(_10567_), .C(_10560_), .Y(_10578_) );
INVX1 INVX1_913 ( .A(decoded_imm_uj_23_), .Y(_10579_) );
INVX1 INVX1_914 ( .A(reg_next_pc_23_), .Y(_10580_) );
NOR2X1 NOR2X1_962 ( .A(_10580_), .B(_10118__bF_buf4), .Y(_10581_) );
AOI21X1 AOI21X1_768 ( .A(_10118__bF_buf3), .B(_4830_), .C(_10581_), .Y(_10582_) );
XNOR2X1 XNOR2X1_35 ( .A(_10582_), .B(_10579_), .Y(_10583_) );
AND2X2 AND2X2_175 ( .A(_10578_), .B(_10583_), .Y(_10584_) );
OAI21X1 OAI21X1_2326 ( .A(_10578_), .B(_10583_), .C(instr_jal_bF_buf5), .Y(_10585_) );
INVX1 INVX1_915 ( .A(_10581_), .Y(_10586_) );
OAI21X1 OAI21X1_2327 ( .A(_4831_), .B(_10103__bF_buf2), .C(_10586_), .Y(_10587_) );
NAND2X1 NAND2X1_708 ( .A(_10561_), .B(_10571_), .Y(_10588_) );
XNOR2X1 XNOR2X1_36 ( .A(_10588_), .B(_10587_), .Y(_10589_) );
OAI21X1 OAI21X1_2328 ( .A(_10589_), .B(_4605__bF_buf1), .C(_10108_), .Y(_10590_) );
OAI21X1 OAI21X1_2329 ( .A(_10584_), .B(_10585_), .C(_10590_), .Y(_10591_) );
NOR2X1 NOR2X1_963 ( .A(_4431__bF_buf2), .B(_10582_), .Y(_10592_) );
OAI21X1 OAI21X1_2330 ( .A(_10099__bF_buf3), .B(_10592_), .C(_10591_), .Y(_10593_) );
AOI21X1 AOI21X1_769 ( .A(_10577_), .B(_10593_), .C(_4426__bF_buf3), .Y(_80__23_) );
NAND2X1 NAND2X1_709 ( .A(reg_next_pc_24_), .B(_4431__bF_buf1), .Y(_10594_) );
INVX1 INVX1_916 ( .A(_4837_), .Y(_10595_) );
OAI21X1 OAI21X1_2331 ( .A(_10109__bF_buf1), .B(_4639__bF_buf3), .C(reg_next_pc_24_), .Y(_10596_) );
OAI21X1 OAI21X1_2332 ( .A(_10595_), .B(_10103__bF_buf1), .C(_10596_), .Y(_10597_) );
NAND2X1 NAND2X1_710 ( .A(cpu_state_1_bF_buf0_), .B(_10597_), .Y(_10598_) );
OAI21X1 OAI21X1_2333 ( .A(_4431__bF_buf0), .B(_4605__bF_buf0), .C(_10598_), .Y(_10599_) );
INVX1 INVX1_917 ( .A(_10583_), .Y(_10600_) );
NAND2X1 NAND2X1_711 ( .A(_10600_), .B(_10563_), .Y(_10601_) );
NOR2X1 NOR2X1_964 ( .A(_10601_), .B(_10566_), .Y(_10602_) );
NAND2X1 NAND2X1_712 ( .A(_10515_), .B(_10602_), .Y(_10603_) );
AOI21X1 AOI21X1_770 ( .A(_10428_), .B(_10421_), .C(_10603_), .Y(_10604_) );
NOR2X1 NOR2X1_965 ( .A(_10579_), .B(_10582_), .Y(_10605_) );
AOI21X1 AOI21X1_771 ( .A(_10560_), .B(_10600_), .C(_10605_), .Y(_10606_) );
OAI21X1 OAI21X1_2334 ( .A(_10565_), .B(_10601_), .C(_10606_), .Y(_10607_) );
AOI21X1 AOI21X1_772 ( .A(_10513_), .B(_10602_), .C(_10607_), .Y(_10608_) );
INVX1 INVX1_918 ( .A(_10608_), .Y(_10609_) );
NOR2X1 NOR2X1_966 ( .A(_10609_), .B(_10604_), .Y(_10610_) );
NAND2X1 NAND2X1_713 ( .A(decoded_imm_uj_24_), .B(_10597_), .Y(_10611_) );
INVX1 INVX1_919 ( .A(decoded_imm_uj_24_), .Y(_10612_) );
INVX1 INVX1_920 ( .A(_10597_), .Y(_10613_) );
NAND2X1 NAND2X1_714 ( .A(_10612_), .B(_10613_), .Y(_10614_) );
NAND2X1 NAND2X1_715 ( .A(_10611_), .B(_10614_), .Y(_10615_) );
OAI21X1 OAI21X1_2335 ( .A(_10610_), .B(_10615_), .C(instr_jal_bF_buf4), .Y(_10616_) );
AOI21X1 AOI21X1_773 ( .A(_10610_), .B(_10615_), .C(_10616_), .Y(_10617_) );
NAND3X1 NAND3X1_64 ( .A(_10561_), .B(_10587_), .C(_10570_), .Y(_10618_) );
NOR2X1 NOR2X1_967 ( .A(_10529_), .B(_10618_), .Y(_10619_) );
NAND2X1 NAND2X1_716 ( .A(_10619_), .B(_10527_), .Y(_10620_) );
XNOR2X1 XNOR2X1_37 ( .A(_10620_), .B(_10613_), .Y(_10621_) );
OAI21X1 OAI21X1_2336 ( .A(_10621_), .B(instr_jal_bF_buf3), .C(decoder_trigger_bF_buf3), .Y(_10622_) );
OAI21X1 OAI21X1_2337 ( .A(_10617_), .B(_10622_), .C(_10599_), .Y(_10623_) );
AOI21X1 AOI21X1_774 ( .A(_10594_), .B(_10623_), .C(_4426__bF_buf2), .Y(_80__24_) );
NAND2X1 NAND2X1_717 ( .A(reg_next_pc_25_), .B(_4431__bF_buf7), .Y(_10624_) );
INVX1 INVX1_921 ( .A(_4849_), .Y(_10625_) );
OAI21X1 OAI21X1_2338 ( .A(_10109__bF_buf0), .B(_4639__bF_buf2), .C(reg_next_pc_25_), .Y(_10626_) );
OAI21X1 OAI21X1_2339 ( .A(_10625_), .B(_10103__bF_buf0), .C(_10626_), .Y(_10627_) );
INVX1 INVX1_922 ( .A(_10627_), .Y(_10628_) );
OAI21X1 OAI21X1_2340 ( .A(_10628_), .B(_4431__bF_buf6), .C(_10123__bF_buf0), .Y(_10629_) );
OAI21X1 OAI21X1_2341 ( .A(_10610_), .B(_10615_), .C(_10611_), .Y(_10630_) );
NAND2X1 NAND2X1_718 ( .A(decoded_imm_uj_25_), .B(_10627_), .Y(_10631_) );
INVX1 INVX1_923 ( .A(decoded_imm_uj_25_), .Y(_10632_) );
NAND2X1 NAND2X1_719 ( .A(_10632_), .B(_10628_), .Y(_10633_) );
NAND2X1 NAND2X1_720 ( .A(_10631_), .B(_10633_), .Y(_10634_) );
INVX1 INVX1_924 ( .A(_10634_), .Y(_10635_) );
OAI21X1 OAI21X1_2342 ( .A(_10630_), .B(_10635_), .C(instr_jal_bF_buf2), .Y(_10636_) );
AOI21X1 AOI21X1_775 ( .A(_10630_), .B(_10635_), .C(_10636_), .Y(_10637_) );
NOR2X1 NOR2X1_968 ( .A(_10613_), .B(_10620_), .Y(_10638_) );
XNOR2X1 XNOR2X1_38 ( .A(_10638_), .B(_10627_), .Y(_10639_) );
OAI21X1 OAI21X1_2343 ( .A(_10639_), .B(instr_jal_bF_buf1), .C(decoder_trigger_bF_buf2), .Y(_10640_) );
OAI21X1 OAI21X1_2344 ( .A(_10637_), .B(_10640_), .C(_10629_), .Y(_10641_) );
AOI21X1 AOI21X1_776 ( .A(_10624_), .B(_10641_), .C(_4426__bF_buf1), .Y(_80__25_) );
NAND2X1 NAND2X1_721 ( .A(reg_next_pc_26_), .B(_4431__bF_buf5), .Y(_10642_) );
INVX1 INVX1_925 ( .A(_4858_), .Y(_10643_) );
OAI21X1 OAI21X1_2345 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_26_), .Y(_10644_) );
OAI21X1 OAI21X1_2346 ( .A(_10643_), .B(_10103__bF_buf6), .C(_10644_), .Y(_10645_) );
NAND2X1 NAND2X1_722 ( .A(cpu_state_1_bF_buf5_), .B(_10645_), .Y(_10646_) );
OAI21X1 OAI21X1_2347 ( .A(_4431__bF_buf4), .B(_4605__bF_buf5), .C(_10646_), .Y(_10647_) );
OAI21X1 OAI21X1_2348 ( .A(_10628_), .B(_10632_), .C(_10611_), .Y(_10648_) );
OAI21X1 OAI21X1_2349 ( .A(decoded_imm_uj_25_), .B(_10627_), .C(_10648_), .Y(_10649_) );
OR2X2 OR2X2_29 ( .A(_10615_), .B(_10634_), .Y(_10650_) );
OAI21X1 OAI21X1_2350 ( .A(_10610_), .B(_10650_), .C(_10649_), .Y(_10651_) );
INVX1 INVX1_926 ( .A(decoded_imm_uj_26_), .Y(_10652_) );
INVX1 INVX1_927 ( .A(_10645_), .Y(_10653_) );
NOR2X1 NOR2X1_969 ( .A(_10652_), .B(_10653_), .Y(_10654_) );
INVX1 INVX1_928 ( .A(_10654_), .Y(_10655_) );
NAND2X1 NAND2X1_723 ( .A(_10652_), .B(_10653_), .Y(_10656_) );
NAND2X1 NAND2X1_724 ( .A(_10656_), .B(_10655_), .Y(_10657_) );
INVX1 INVX1_929 ( .A(_10657_), .Y(_10658_) );
OAI21X1 OAI21X1_2351 ( .A(_10651_), .B(_10658_), .C(instr_jal_bF_buf0), .Y(_10659_) );
AOI21X1 AOI21X1_777 ( .A(_10651_), .B(_10658_), .C(_10659_), .Y(_10660_) );
OR2X2 OR2X2_30 ( .A(_10618_), .B(_10492_), .Y(_10661_) );
NOR2X1 NOR2X1_970 ( .A(_10628_), .B(_10613_), .Y(_10662_) );
INVX1 INVX1_930 ( .A(_10662_), .Y(_10663_) );
NOR3X1 NOR3X1_3 ( .A(_10661_), .B(_10663_), .C(_10482_), .Y(_10664_) );
XNOR2X1 XNOR2X1_39 ( .A(_10664_), .B(_10645_), .Y(_10665_) );
OAI21X1 OAI21X1_2352 ( .A(_10665_), .B(instr_jal_bF_buf6), .C(decoder_trigger_bF_buf1), .Y(_10666_) );
OAI21X1 OAI21X1_2353 ( .A(_10660_), .B(_10666_), .C(_10647_), .Y(_10667_) );
AOI21X1 AOI21X1_778 ( .A(_10642_), .B(_10667_), .C(_4426__bF_buf0), .Y(_80__26_) );
NAND2X1 NAND2X1_725 ( .A(reg_next_pc_27_), .B(_4431__bF_buf3), .Y(_10668_) );
AOI21X1 AOI21X1_779 ( .A(_10658_), .B(_10651_), .C(_10654_), .Y(_10669_) );
INVX1 INVX1_931 ( .A(decoded_imm_uj_27_), .Y(_10670_) );
OAI21X1 OAI21X1_2354 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_27_), .Y(_10671_) );
OAI21X1 OAI21X1_2355 ( .A(_4869_), .B(_10103__bF_buf5), .C(_10671_), .Y(_10672_) );
INVX1 INVX1_932 ( .A(_10672_), .Y(_10673_) );
XNOR2X1 XNOR2X1_40 ( .A(_10673_), .B(_10670_), .Y(_10674_) );
AND2X2 AND2X2_176 ( .A(_10669_), .B(_10674_), .Y(_10675_) );
OAI21X1 OAI21X1_2356 ( .A(_10669_), .B(_10674_), .C(instr_jal_bF_buf5), .Y(_10676_) );
NAND3X1 NAND3X1_65 ( .A(_10645_), .B(_10672_), .C(_10664_), .Y(_10677_) );
NAND2X1 NAND2X1_726 ( .A(_10645_), .B(_10664_), .Y(_10678_) );
AOI21X1 AOI21X1_780 ( .A(_10673_), .B(_10678_), .C(instr_jal_bF_buf4), .Y(_10679_) );
AOI21X1 AOI21X1_781 ( .A(_10677_), .B(_10679_), .C(_4605__bF_buf4), .Y(_10680_) );
OAI21X1 OAI21X1_2357 ( .A(_10675_), .B(_10676_), .C(_10680_), .Y(_10681_) );
NOR2X1 NOR2X1_971 ( .A(_4431__bF_buf2), .B(_10673_), .Y(_10682_) );
OAI21X1 OAI21X1_2358 ( .A(_10099__bF_buf2), .B(_10682_), .C(_10681_), .Y(_10683_) );
AOI21X1 AOI21X1_782 ( .A(_10668_), .B(_10683_), .C(_4426__bF_buf11), .Y(_80__27_) );
NAND2X1 NAND2X1_727 ( .A(reg_next_pc_28_), .B(_4431__bF_buf1), .Y(_10684_) );
INVX1 INVX1_933 ( .A(_4875_), .Y(_10685_) );
OAI21X1 OAI21X1_2359 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_28_), .Y(_10686_) );
OAI21X1 OAI21X1_2360 ( .A(_10685_), .B(_10103__bF_buf4), .C(_10686_), .Y(_10687_) );
NAND2X1 NAND2X1_728 ( .A(cpu_state_1_bF_buf4_), .B(_10687_), .Y(_10688_) );
OAI21X1 OAI21X1_2361 ( .A(_4431__bF_buf0), .B(_4605__bF_buf3), .C(_10688_), .Y(_10689_) );
INVX1 INVX1_934 ( .A(_10687_), .Y(_10690_) );
OAI21X1 OAI21X1_2362 ( .A(_10677_), .B(_10690_), .C(_4499__bF_buf3), .Y(_10691_) );
AOI21X1 AOI21X1_783 ( .A(_10677_), .B(_10690_), .C(_10691_), .Y(_10692_) );
OR2X2 OR2X2_31 ( .A(_10657_), .B(_10674_), .Y(_10693_) );
OR2X2 OR2X2_32 ( .A(_10693_), .B(_10650_), .Y(_10694_) );
NOR2X1 NOR2X1_972 ( .A(_10649_), .B(_10693_), .Y(_10695_) );
OAI21X1 OAI21X1_2363 ( .A(decoded_imm_uj_27_), .B(_10672_), .C(_10654_), .Y(_10696_) );
OAI21X1 OAI21X1_2364 ( .A(_10670_), .B(_10673_), .C(_10696_), .Y(_10697_) );
NOR2X1 NOR2X1_973 ( .A(_10697_), .B(_10695_), .Y(_10698_) );
OAI21X1 OAI21X1_2365 ( .A(_10610_), .B(_10694_), .C(_10698_), .Y(_10699_) );
INVX1 INVX1_935 ( .A(decoded_imm_uj_28_), .Y(_10700_) );
NAND2X1 NAND2X1_729 ( .A(_10700_), .B(_10690_), .Y(_10701_) );
NOR2X1 NOR2X1_974 ( .A(_10700_), .B(_10690_), .Y(_10702_) );
INVX1 INVX1_936 ( .A(_10702_), .Y(_10703_) );
NAND2X1 NAND2X1_730 ( .A(_10701_), .B(_10703_), .Y(_10704_) );
INVX1 INVX1_937 ( .A(_10704_), .Y(_10705_) );
XNOR2X1 XNOR2X1_41 ( .A(_10699_), .B(_10705_), .Y(_10706_) );
OAI21X1 OAI21X1_2366 ( .A(_10706_), .B(_4499__bF_buf2), .C(decoder_trigger_bF_buf0), .Y(_10707_) );
OAI21X1 OAI21X1_2367 ( .A(_10707_), .B(_10692_), .C(_10689_), .Y(_10708_) );
AOI21X1 AOI21X1_784 ( .A(_10684_), .B(_10708_), .C(_4426__bF_buf10), .Y(_80__28_) );
NAND2X1 NAND2X1_731 ( .A(reg_next_pc_29_), .B(_4431__bF_buf7), .Y(_10709_) );
AOI21X1 AOI21X1_785 ( .A(_10705_), .B(_10699_), .C(_10702_), .Y(_10710_) );
OAI21X1 OAI21X1_2368 ( .A(_10109__bF_buf1), .B(_4639__bF_buf3), .C(reg_next_pc_29_), .Y(_10711_) );
INVX1 INVX1_938 ( .A(_10711_), .Y(_10712_) );
AOI21X1 AOI21X1_786 ( .A(_10118__bF_buf2), .B(_4888_), .C(_10712_), .Y(_10713_) );
INVX1 INVX1_939 ( .A(_10713_), .Y(_10714_) );
NOR2X1 NOR2X1_975 ( .A(decoded_imm_uj_29_), .B(_10714_), .Y(_10715_) );
INVX1 INVX1_940 ( .A(decoded_imm_uj_29_), .Y(_10716_) );
NOR2X1 NOR2X1_976 ( .A(_10716_), .B(_10713_), .Y(_10717_) );
NOR2X1 NOR2X1_977 ( .A(_10717_), .B(_10715_), .Y(_10718_) );
INVX1 INVX1_941 ( .A(_10718_), .Y(_10719_) );
AND2X2 AND2X2_177 ( .A(_10710_), .B(_10719_), .Y(_10720_) );
OAI21X1 OAI21X1_2369 ( .A(_10710_), .B(_10719_), .C(instr_jal_bF_buf3), .Y(_10721_) );
NAND3X1 NAND3X1_66 ( .A(_10645_), .B(_10672_), .C(_10662_), .Y(_10722_) );
NOR2X1 NOR2X1_978 ( .A(_10722_), .B(_10620_), .Y(_10723_) );
NAND2X1 NAND2X1_732 ( .A(_10687_), .B(_10723_), .Y(_1120_) );
XNOR2X1 XNOR2X1_42 ( .A(_1120_), .B(_10714_), .Y(_1121_) );
OAI21X1 OAI21X1_2370 ( .A(_1121_), .B(_4605__bF_buf2), .C(_10108_), .Y(_1122_) );
OAI21X1 OAI21X1_2371 ( .A(_10720_), .B(_10721_), .C(_1122_), .Y(_1123_) );
NOR2X1 NOR2X1_979 ( .A(_4431__bF_buf6), .B(_10713_), .Y(_1124_) );
OAI21X1 OAI21X1_2372 ( .A(_10099__bF_buf1), .B(_1124_), .C(_1123_), .Y(_1125_) );
AOI21X1 AOI21X1_787 ( .A(_10709_), .B(_1125_), .C(_4426__bF_buf9), .Y(_80__29_) );
NAND2X1 NAND2X1_733 ( .A(reg_next_pc_30_), .B(_4431__bF_buf5), .Y(_1126_) );
INVX1 INVX1_942 ( .A(_4897_), .Y(_1127_) );
OAI21X1 OAI21X1_2373 ( .A(_10109__bF_buf0), .B(_4639__bF_buf2), .C(reg_next_pc_30_), .Y(_1128_) );
OAI21X1 OAI21X1_2374 ( .A(_1127_), .B(_10103__bF_buf3), .C(_1128_), .Y(_1129_) );
NAND2X1 NAND2X1_734 ( .A(cpu_state_1_bF_buf3_), .B(_1129_), .Y(_1130_) );
OAI21X1 OAI21X1_2375 ( .A(_4431__bF_buf4), .B(_4605__bF_buf1), .C(_1130_), .Y(_1131_) );
NOR3X1 NOR3X1_4 ( .A(_10690_), .B(_10713_), .C(_10677_), .Y(_1132_) );
OAI21X1 OAI21X1_2376 ( .A(_1132_), .B(_1129_), .C(_4499__bF_buf1), .Y(_1133_) );
AOI21X1 AOI21X1_788 ( .A(_1132_), .B(_1129_), .C(_1133_), .Y(_1134_) );
NOR2X1 NOR2X1_980 ( .A(_10650_), .B(_10693_), .Y(_1135_) );
OAI21X1 OAI21X1_2377 ( .A(_10604_), .B(_10609_), .C(_1135_), .Y(_1136_) );
NOR2X1 NOR2X1_981 ( .A(_10704_), .B(_10719_), .Y(_1137_) );
INVX1 INVX1_943 ( .A(_1137_), .Y(_1138_) );
AOI21X1 AOI21X1_789 ( .A(_10698_), .B(_1136_), .C(_1138_), .Y(_1139_) );
AOI21X1 AOI21X1_790 ( .A(_10702_), .B(_10718_), .C(_10717_), .Y(_1140_) );
INVX1 INVX1_944 ( .A(_1140_), .Y(_1141_) );
NOR2X1 NOR2X1_982 ( .A(_1141_), .B(_1139_), .Y(_1142_) );
NOR2X1 NOR2X1_983 ( .A(decoded_imm_uj_30_), .B(_1129_), .Y(_1143_) );
NAND2X1 NAND2X1_735 ( .A(decoded_imm_uj_30_), .B(_1129_), .Y(_1144_) );
INVX1 INVX1_945 ( .A(_1144_), .Y(_1145_) );
NOR2X1 NOR2X1_984 ( .A(_1143_), .B(_1145_), .Y(_1146_) );
INVX1 INVX1_946 ( .A(_1146_), .Y(_1147_) );
AND2X2 AND2X2_178 ( .A(_1142_), .B(_1147_), .Y(_1148_) );
OAI21X1 OAI21X1_2378 ( .A(_1142_), .B(_1147_), .C(instr_jal_bF_buf2), .Y(_1149_) );
OAI21X1 OAI21X1_2379 ( .A(_1148_), .B(_1149_), .C(decoder_trigger_bF_buf3), .Y(_1150_) );
OAI21X1 OAI21X1_2380 ( .A(_1150_), .B(_1134_), .C(_1131_), .Y(_1151_) );
AOI21X1 AOI21X1_791 ( .A(_1126_), .B(_1151_), .C(_4426__bF_buf8), .Y(_80__30_) );
NAND2X1 NAND2X1_736 ( .A(reg_next_pc_31_), .B(_4431__bF_buf3), .Y(_1152_) );
NAND2X1 NAND2X1_737 ( .A(_10150_), .B(_10143_), .Y(_1153_) );
NAND2X1 NAND2X1_738 ( .A(_10168_), .B(_1153_), .Y(_1154_) );
NOR3X1 NOR3X1_5 ( .A(_10136_), .B(_1154_), .C(_10128_), .Y(_1155_) );
NOR2X1 NOR2X1_985 ( .A(_10209_), .B(_10255_), .Y(_1156_) );
OAI21X1 OAI21X1_2381 ( .A(_1155_), .B(_10169_), .C(_1156_), .Y(_1157_) );
AOI21X1 AOI21X1_792 ( .A(_10294_), .B(_1157_), .C(_10438_), .Y(_1158_) );
INVX1 INVX1_947 ( .A(_10428_), .Y(_1159_) );
OR2X2 OR2X2_33 ( .A(_10511_), .B(_10514_), .Y(_1160_) );
NOR3X1 NOR3X1_6 ( .A(_10560_), .B(_10562_), .C(_10583_), .Y(_1161_) );
NAND3X1 NAND3X1_67 ( .A(_10521_), .B(_10545_), .C(_1161_), .Y(_1162_) );
NOR2X1 NOR2X1_986 ( .A(_1162_), .B(_1160_), .Y(_1163_) );
OAI21X1 OAI21X1_2382 ( .A(_1158_), .B(_1159_), .C(_1163_), .Y(_1164_) );
AOI21X1 AOI21X1_793 ( .A(_10608_), .B(_1164_), .C(_10694_), .Y(_1165_) );
OR2X2 OR2X2_34 ( .A(_10695_), .B(_10697_), .Y(_1166_) );
OAI21X1 OAI21X1_2383 ( .A(_1165_), .B(_1166_), .C(_1137_), .Y(_1167_) );
AOI21X1 AOI21X1_794 ( .A(_1140_), .B(_1167_), .C(_1147_), .Y(_1168_) );
INVX1 INVX1_948 ( .A(decoded_imm_uj_31_), .Y(_1169_) );
OAI21X1 OAI21X1_2384 ( .A(_10109__bF_buf4), .B(_4639__bF_buf1), .C(reg_next_pc_31_), .Y(_1170_) );
INVX1 INVX1_949 ( .A(_1170_), .Y(_1171_) );
AOI21X1 AOI21X1_795 ( .A(_10118__bF_buf1), .B(_4905_), .C(_1171_), .Y(_1172_) );
XNOR2X1 XNOR2X1_43 ( .A(_1172_), .B(_1169_), .Y(_1173_) );
OAI21X1 OAI21X1_2385 ( .A(_1168_), .B(_1145_), .C(_1173_), .Y(_1174_) );
OAI21X1 OAI21X1_2386 ( .A(_1139_), .B(_1141_), .C(_1146_), .Y(_1175_) );
INVX1 INVX1_950 ( .A(_1173_), .Y(_1176_) );
NAND3X1 NAND3X1_68 ( .A(_1144_), .B(_1176_), .C(_1175_), .Y(_1177_) );
AOI21X1 AOI21X1_796 ( .A(_1177_), .B(_1174_), .C(_4499__bF_buf0), .Y(_1178_) );
NAND3X1 NAND3X1_69 ( .A(_1129_), .B(_1172_), .C(_1132_), .Y(_1179_) );
INVX1 INVX1_951 ( .A(_1172_), .Y(_1180_) );
NOR2X1 NOR2X1_987 ( .A(_10713_), .B(_10690_), .Y(_1181_) );
NAND3X1 NAND3X1_70 ( .A(_1129_), .B(_1181_), .C(_10723_), .Y(_1182_) );
AOI21X1 AOI21X1_797 ( .A(_1180_), .B(_1182_), .C(_4605__bF_buf0), .Y(_1183_) );
AOI21X1 AOI21X1_798 ( .A(_1183_), .B(_1179_), .C(_10107_), .Y(_1184_) );
OAI21X1 OAI21X1_2387 ( .A(_1172_), .B(_4431__bF_buf2), .C(_10123__bF_buf4), .Y(_1185_) );
OAI21X1 OAI21X1_2388 ( .A(_1178_), .B(_1184_), .C(_1185_), .Y(_1186_) );
AOI21X1 AOI21X1_799 ( .A(_1152_), .B(_1186_), .C(_4426__bF_buf7), .Y(_80__31_) );
OAI21X1 OAI21X1_2389 ( .A(cpu_state_1_bF_buf2_), .B(reg_pc_0_), .C(resetn_bF_buf11), .Y(_1187_) );
AOI21X1 AOI21X1_800 ( .A(cpu_state_1_bF_buf1_), .B(_10110_), .C(_1187_), .Y(_84__0_) );
NAND2X1 NAND2X1_739 ( .A(reg_pc_1_), .B(_4431__bF_buf1), .Y(_1188_) );
AOI21X1 AOI21X1_801 ( .A(_1188_), .B(_10124_), .C(_4426__bF_buf6), .Y(_84__1_) );
OAI21X1 OAI21X1_2390 ( .A(cpu_state_1_bF_buf0_), .B(reg_pc_2_), .C(resetn_bF_buf10), .Y(_1189_) );
AOI21X1 AOI21X1_802 ( .A(cpu_state_1_bF_buf5_), .B(_10134_), .C(_1189_), .Y(_84__2_) );
AOI21X1 AOI21X1_803 ( .A(_4431__bF_buf0), .B(reg_pc_3_), .C(_10144_), .Y(_1190_) );
NOR2X1 NOR2X1_988 ( .A(_4426__bF_buf5), .B(_1190_), .Y(_84__3_) );
MUX2X1 MUX2X1_217 ( .A(_10166_), .B(reg_pc_4_), .S(cpu_state_1_bF_buf4_), .Y(_1191_) );
NOR2X1 NOR2X1_989 ( .A(_4426__bF_buf4), .B(_1191_), .Y(_84__4_) );
MUX2X1 MUX2X1_218 ( .A(_10192_), .B(reg_pc_5_), .S(cpu_state_1_bF_buf3_), .Y(_1192_) );
NOR2X1 NOR2X1_990 ( .A(_4426__bF_buf3), .B(_1192_), .Y(_84__5_) );
MUX2X1 MUX2X1_219 ( .A(_10206_), .B(reg_pc_6_), .S(cpu_state_1_bF_buf2_), .Y(_1193_) );
NOR2X1 NOR2X1_991 ( .A(_4426__bF_buf2), .B(_1193_), .Y(_84__6_) );
MUX2X1 MUX2X1_220 ( .A(_10227_), .B(reg_pc_7_), .S(cpu_state_1_bF_buf1_), .Y(_1194_) );
NOR2X1 NOR2X1_992 ( .A(_4426__bF_buf1), .B(_1194_), .Y(_84__7_) );
AOI21X1 AOI21X1_804 ( .A(_4431__bF_buf7), .B(reg_pc_8_), .C(_10243_), .Y(_1195_) );
NOR2X1 NOR2X1_993 ( .A(_4426__bF_buf0), .B(_1195_), .Y(_84__8_) );
MUX2X1 MUX2X1_221 ( .A(_10272_), .B(reg_pc_9_), .S(cpu_state_1_bF_buf0_), .Y(_1196_) );
NOR2X1 NOR2X1_994 ( .A(_4426__bF_buf11), .B(_1196_), .Y(_84__9_) );
MUX2X1 MUX2X1_222 ( .A(_10285_), .B(reg_pc_10_), .S(cpu_state_1_bF_buf5_), .Y(_1197_) );
NOR2X1 NOR2X1_995 ( .A(_4426__bF_buf10), .B(_1197_), .Y(_84__10_) );
AOI21X1 AOI21X1_805 ( .A(_4431__bF_buf6), .B(reg_pc_11_), .C(_10327_), .Y(_1198_) );
NOR2X1 NOR2X1_996 ( .A(_4426__bF_buf9), .B(_1198_), .Y(_84__11_) );
OAI21X1 OAI21X1_2391 ( .A(cpu_state_1_bF_buf4_), .B(_4719_), .C(_10332_), .Y(_1199_) );
AND2X2 AND2X2_179 ( .A(_1199_), .B(resetn_bF_buf9), .Y(_84__12_) );
AOI21X1 AOI21X1_806 ( .A(_4431__bF_buf5), .B(reg_pc_13_), .C(_10375_), .Y(_1200_) );
NOR2X1 NOR2X1_997 ( .A(_4426__bF_buf8), .B(_1200_), .Y(_84__13_) );
MUX2X1 MUX2X1_223 ( .A(_10379_), .B(reg_pc_14_), .S(cpu_state_1_bF_buf3_), .Y(_1201_) );
NOR2X1 NOR2X1_998 ( .A(_4426__bF_buf7), .B(_1201_), .Y(_84__14_) );
MUX2X1 MUX2X1_224 ( .A(_10399_), .B(reg_pc_15_), .S(cpu_state_1_bF_buf2_), .Y(_1202_) );
NOR2X1 NOR2X1_999 ( .A(_4426__bF_buf6), .B(_1202_), .Y(_84__15_) );
MUX2X1 MUX2X1_225 ( .A(_10431_), .B(reg_pc_16_), .S(cpu_state_1_bF_buf1_), .Y(_1203_) );
NOR2X1 NOR2X1_1000 ( .A(_4426__bF_buf5), .B(_1203_), .Y(_84__16_) );
AOI21X1 AOI21X1_807 ( .A(_4431__bF_buf4), .B(reg_pc_17_), .C(_10465_), .Y(_1204_) );
NOR2X1 NOR2X1_1001 ( .A(_4426__bF_buf4), .B(_1204_), .Y(_84__17_) );
MUX2X1 MUX2X1_226 ( .A(_10474_), .B(reg_pc_18_), .S(cpu_state_1_bF_buf0_), .Y(_1205_) );
NOR2X1 NOR2X1_1002 ( .A(_4426__bF_buf3), .B(_1205_), .Y(_84__18_) );
MUX2X1 MUX2X1_227 ( .A(_10495_), .B(reg_pc_19_), .S(cpu_state_1_bF_buf5_), .Y(_1206_) );
NOR2X1 NOR2X1_1003 ( .A(_4426__bF_buf2), .B(_1206_), .Y(_84__19_) );
AOI21X1 AOI21X1_808 ( .A(_4431__bF_buf3), .B(reg_pc_20_), .C(_10509_), .Y(_1207_) );
NOR2X1 NOR2X1_1004 ( .A(_4426__bF_buf1), .B(_1207_), .Y(_84__20_) );
MUX2X1 MUX2X1_228 ( .A(_10543_), .B(reg_pc_21_), .S(cpu_state_1_bF_buf4_), .Y(_1208_) );
NOR2X1 NOR2X1_1005 ( .A(_4426__bF_buf0), .B(_1208_), .Y(_84__21_) );
MUX2X1 MUX2X1_229 ( .A(_10561_), .B(reg_pc_22_), .S(cpu_state_1_bF_buf3_), .Y(_1209_) );
NOR2X1 NOR2X1_1006 ( .A(_4426__bF_buf11), .B(_1209_), .Y(_84__22_) );
AOI21X1 AOI21X1_809 ( .A(_4431__bF_buf2), .B(reg_pc_23_), .C(_10592_), .Y(_1210_) );
NOR2X1 NOR2X1_1007 ( .A(_4426__bF_buf10), .B(_1210_), .Y(_84__23_) );
OAI21X1 OAI21X1_2392 ( .A(cpu_state_1_bF_buf2_), .B(_4841_), .C(_10598_), .Y(_1211_) );
AND2X2 AND2X2_180 ( .A(_1211_), .B(resetn_bF_buf8), .Y(_84__24_) );
MUX2X1 MUX2X1_230 ( .A(_10627_), .B(reg_pc_25_), .S(cpu_state_1_bF_buf1_), .Y(_1212_) );
NOR2X1 NOR2X1_1008 ( .A(_4426__bF_buf9), .B(_1212_), .Y(_84__25_) );
OAI21X1 OAI21X1_2393 ( .A(cpu_state_1_bF_buf0_), .B(_4860_), .C(_10646_), .Y(_1213_) );
AND2X2 AND2X2_181 ( .A(_1213_), .B(resetn_bF_buf7), .Y(_84__26_) );
AOI21X1 AOI21X1_810 ( .A(_4431__bF_buf1), .B(reg_pc_27_), .C(_10682_), .Y(_1214_) );
NOR2X1 NOR2X1_1009 ( .A(_4426__bF_buf8), .B(_1214_), .Y(_84__27_) );
INVX1 INVX1_952 ( .A(reg_pc_28_), .Y(_1215_) );
OAI21X1 OAI21X1_2394 ( .A(cpu_state_1_bF_buf5_), .B(_1215_), .C(_10688_), .Y(_1216_) );
AND2X2 AND2X2_182 ( .A(_1216_), .B(resetn_bF_buf6), .Y(_84__28_) );
AOI21X1 AOI21X1_811 ( .A(_4431__bF_buf0), .B(reg_pc_29_), .C(_1124_), .Y(_1217_) );
NOR2X1 NOR2X1_1010 ( .A(_4426__bF_buf7), .B(_1217_), .Y(_84__29_) );
OAI21X1 OAI21X1_2395 ( .A(cpu_state_1_bF_buf4_), .B(_4898_), .C(_1130_), .Y(_1218_) );
AND2X2 AND2X2_183 ( .A(_1218_), .B(resetn_bF_buf5), .Y(_84__30_) );
MUX2X1 MUX2X1_231 ( .A(_1180_), .B(reg_pc_31_), .S(cpu_state_1_bF_buf3_), .Y(_1219_) );
NOR2X1 NOR2X1_1011 ( .A(_4426__bF_buf6), .B(_1219_), .Y(_84__31_) );
OAI21X1 OAI21X1_2396 ( .A(_10099__bF_buf0), .B(count_instr_0_), .C(resetn_bF_buf4), .Y(_1220_) );
AOI21X1 AOI21X1_812 ( .A(count_instr_0_), .B(_10099__bF_buf3), .C(_1220_), .Y(_1__0_) );
AOI21X1 AOI21X1_813 ( .A(count_instr_0_), .B(_10099__bF_buf2), .C(count_instr_1_), .Y(_1221_) );
NAND2X1 NAND2X1_740 ( .A(count_instr_0_), .B(count_instr_1_), .Y(_1222_) );
OAI21X1 OAI21X1_2397 ( .A(_10123__bF_buf3), .B(_1222_), .C(resetn_bF_buf3), .Y(_1223_) );
NOR2X1 NOR2X1_1012 ( .A(_1221_), .B(_1223_), .Y(_1__1_) );
NOR2X1 NOR2X1_1013 ( .A(_1222_), .B(_10123__bF_buf2), .Y(_1224_) );
AND2X2 AND2X2_184 ( .A(_1224_), .B(count_instr_2_), .Y(_1225_) );
OAI21X1 OAI21X1_2398 ( .A(_1224_), .B(count_instr_2_), .C(resetn_bF_buf2), .Y(_1226_) );
NOR2X1 NOR2X1_1014 ( .A(_1226_), .B(_1225_), .Y(_1__2_) );
NAND2X1 NAND2X1_741 ( .A(count_instr_2_), .B(count_instr_3_), .Y(_1227_) );
NOR2X1 NOR2X1_1015 ( .A(_1222_), .B(_1227_), .Y(_1228_) );
INVX1 INVX1_953 ( .A(_1228_), .Y(_1229_) );
NOR2X1 NOR2X1_1016 ( .A(_10123__bF_buf1), .B(_1229_), .Y(_1230_) );
OAI21X1 OAI21X1_2399 ( .A(_1225_), .B(count_instr_3_), .C(resetn_bF_buf1), .Y(_1231_) );
NOR2X1 NOR2X1_1017 ( .A(_1230_), .B(_1231_), .Y(_1__3_) );
NAND2X1 NAND2X1_742 ( .A(count_instr_4_), .B(_1230_), .Y(_1232_) );
INVX1 INVX1_954 ( .A(_1232_), .Y(_1233_) );
OAI21X1 OAI21X1_2400 ( .A(_1230_), .B(count_instr_4_), .C(resetn_bF_buf0), .Y(_1234_) );
NOR2X1 NOR2X1_1018 ( .A(_1234_), .B(_1233_), .Y(_1__4_) );
INVX1 INVX1_955 ( .A(count_instr_5_), .Y(_1235_) );
OAI21X1 OAI21X1_2401 ( .A(_1232_), .B(_1235_), .C(resetn_bF_buf11), .Y(_1236_) );
AOI21X1 AOI21X1_814 ( .A(_1235_), .B(_1232_), .C(_1236_), .Y(_1__5_) );
OAI21X1 OAI21X1_2402 ( .A(_1232_), .B(_1235_), .C(count_instr_6_), .Y(_1237_) );
INVX1 INVX1_956 ( .A(count_instr_6_), .Y(_1238_) );
NAND3X1 NAND3X1_71 ( .A(count_instr_5_), .B(_1238_), .C(_1233_), .Y(_1239_) );
AOI21X1 AOI21X1_815 ( .A(_1237_), .B(_1239_), .C(_4426__bF_buf5), .Y(_1__6_) );
NAND2X1 NAND2X1_743 ( .A(count_instr_4_), .B(count_instr_5_), .Y(_1240_) );
NOR2X1 NOR2X1_1019 ( .A(_1240_), .B(_1229_), .Y(_1241_) );
INVX1 INVX1_957 ( .A(_1241_), .Y(_1242_) );
NAND2X1 NAND2X1_744 ( .A(count_instr_6_), .B(count_instr_7_), .Y(_1243_) );
NOR2X1 NOR2X1_1020 ( .A(_1243_), .B(_1242_), .Y(_1244_) );
NAND2X1 NAND2X1_745 ( .A(_10099__bF_buf1), .B(_1244_), .Y(_1245_) );
INVX1 INVX1_958 ( .A(_1245_), .Y(_1246_) );
NAND2X1 NAND2X1_746 ( .A(count_instr_6_), .B(_10099__bF_buf0), .Y(_1247_) );
NOR2X1 NOR2X1_1021 ( .A(_1247_), .B(_1242_), .Y(_1248_) );
OAI21X1 OAI21X1_2403 ( .A(_1248_), .B(count_instr_7_), .C(resetn_bF_buf10), .Y(_1249_) );
NOR2X1 NOR2X1_1022 ( .A(_1249_), .B(_1246_), .Y(_1__7_) );
OAI21X1 OAI21X1_2404 ( .A(_1246_), .B(count_instr_8_), .C(resetn_bF_buf9), .Y(_1250_) );
AOI21X1 AOI21X1_816 ( .A(count_instr_8_), .B(_1246_), .C(_1250_), .Y(_1__8_) );
AOI21X1 AOI21X1_817 ( .A(count_instr_8_), .B(_1246_), .C(count_instr_9_), .Y(_1251_) );
NAND2X1 NAND2X1_747 ( .A(count_instr_8_), .B(count_instr_9_), .Y(_1252_) );
OAI21X1 OAI21X1_2405 ( .A(_1245_), .B(_1252_), .C(resetn_bF_buf8), .Y(_1253_) );
NOR2X1 NOR2X1_1023 ( .A(_1253_), .B(_1251_), .Y(_1__9_) );
NOR2X1 NOR2X1_1024 ( .A(_1252_), .B(_1245_), .Y(_1254_) );
OAI21X1 OAI21X1_2406 ( .A(_1254_), .B(count_instr_10_), .C(resetn_bF_buf7), .Y(_1255_) );
AOI21X1 AOI21X1_818 ( .A(count_instr_10_), .B(_1254_), .C(_1255_), .Y(_1__10_) );
AOI21X1 AOI21X1_819 ( .A(count_instr_10_), .B(_1254_), .C(count_instr_11_), .Y(_1256_) );
NAND2X1 NAND2X1_748 ( .A(count_instr_10_), .B(count_instr_11_), .Y(_1257_) );
INVX1 INVX1_959 ( .A(_1257_), .Y(_1258_) );
NAND2X1 NAND2X1_749 ( .A(_1258_), .B(_1254_), .Y(_1259_) );
NAND2X1 NAND2X1_750 ( .A(resetn_bF_buf6), .B(_1259_), .Y(_1260_) );
NOR2X1 NOR2X1_1025 ( .A(_1256_), .B(_1260_), .Y(_1__11_) );
NAND2X1 NAND2X1_751 ( .A(count_instr_12_), .B(_1259_), .Y(_1261_) );
OR2X2 OR2X2_35 ( .A(_1259_), .B(count_instr_12_), .Y(_1262_) );
AOI21X1 AOI21X1_820 ( .A(_1261_), .B(_1262_), .C(_4426__bF_buf4), .Y(_1__12_) );
NOR2X1 NOR2X1_1026 ( .A(_1240_), .B(_1243_), .Y(_1263_) );
NAND2X1 NAND2X1_752 ( .A(_1228_), .B(_1263_), .Y(_1264_) );
INVX1 INVX1_960 ( .A(_1252_), .Y(_1265_) );
NAND2X1 NAND2X1_753 ( .A(_1265_), .B(_1258_), .Y(_1266_) );
NOR2X1 NOR2X1_1027 ( .A(_1266_), .B(_1264_), .Y(_1267_) );
NAND3X1 NAND3X1_72 ( .A(count_instr_12_), .B(_10099__bF_buf3), .C(_1267_), .Y(_1268_) );
XNOR2X1 XNOR2X1_44 ( .A(_1268_), .B(count_instr_13_), .Y(_1269_) );
AND2X2 AND2X2_185 ( .A(_1269_), .B(resetn_bF_buf5), .Y(_1__13_) );
INVX1 INVX1_961 ( .A(count_instr_13_), .Y(_1270_) );
NOR2X1 NOR2X1_1028 ( .A(_1270_), .B(_1268_), .Y(_1271_) );
XNOR2X1 XNOR2X1_45 ( .A(_1271_), .B(count_instr_14_), .Y(_1272_) );
NOR2X1 NOR2X1_1029 ( .A(_4426__bF_buf3), .B(_1272_), .Y(_1__14_) );
NAND2X1 NAND2X1_754 ( .A(count_instr_12_), .B(_1265_), .Y(_1273_) );
NOR2X1 NOR2X1_1030 ( .A(_1257_), .B(_1273_), .Y(_1274_) );
NAND3X1 NAND3X1_73 ( .A(count_instr_13_), .B(count_instr_14_), .C(_1274_), .Y(_1275_) );
NOR2X1 NOR2X1_1031 ( .A(_1275_), .B(_1245_), .Y(_1276_) );
OAI21X1 OAI21X1_2407 ( .A(_1276_), .B(count_instr_15_), .C(resetn_bF_buf4), .Y(_1277_) );
AOI21X1 AOI21X1_821 ( .A(count_instr_15_), .B(_1276_), .C(_1277_), .Y(_1__15_) );
INVX1 INVX1_962 ( .A(count_instr_16_), .Y(_1278_) );
NAND2X1 NAND2X1_755 ( .A(count_instr_15_), .B(_1276_), .Y(_1279_) );
XNOR2X1 XNOR2X1_46 ( .A(_1279_), .B(_1278_), .Y(_1280_) );
NOR2X1 NOR2X1_1032 ( .A(_4426__bF_buf2), .B(_1280_), .Y(_1__16_) );
NAND2X1 NAND2X1_756 ( .A(count_instr_12_), .B(count_instr_13_), .Y(_1281_) );
NAND2X1 NAND2X1_757 ( .A(count_instr_14_), .B(count_instr_15_), .Y(_1282_) );
NOR2X1 NOR2X1_1033 ( .A(_1281_), .B(_1282_), .Y(_1283_) );
NAND3X1 NAND3X1_74 ( .A(_1265_), .B(_1258_), .C(_1283_), .Y(_1284_) );
NOR2X1 NOR2X1_1034 ( .A(_1264_), .B(_1284_), .Y(_1285_) );
INVX1 INVX1_963 ( .A(_1285_), .Y(_1286_) );
NAND2X1 NAND2X1_758 ( .A(count_instr_16_), .B(_10099__bF_buf2), .Y(_1287_) );
NOR2X1 NOR2X1_1035 ( .A(_1287_), .B(_1286_), .Y(_1288_) );
NAND2X1 NAND2X1_759 ( .A(count_instr_17_), .B(_1288_), .Y(_1289_) );
INVX1 INVX1_964 ( .A(_1289_), .Y(_1290_) );
OAI21X1 OAI21X1_2408 ( .A(_1288_), .B(count_instr_17_), .C(resetn_bF_buf3), .Y(_1291_) );
NOR2X1 NOR2X1_1036 ( .A(_1291_), .B(_1290_), .Y(_1__17_) );
NAND2X1 NAND2X1_760 ( .A(count_instr_18_), .B(_1289_), .Y(_1292_) );
OR2X2 OR2X2_36 ( .A(_1289_), .B(count_instr_18_), .Y(_1293_) );
AOI21X1 AOI21X1_822 ( .A(_1292_), .B(_1293_), .C(_4426__bF_buf1), .Y(_1__18_) );
INVX1 INVX1_965 ( .A(count_instr_19_), .Y(_1294_) );
NAND2X1 NAND2X1_761 ( .A(count_instr_18_), .B(_1290_), .Y(_1295_) );
OAI21X1 OAI21X1_2409 ( .A(_1295_), .B(_1294_), .C(resetn_bF_buf2), .Y(_1296_) );
AOI21X1 AOI21X1_823 ( .A(_1294_), .B(_1295_), .C(_1296_), .Y(_1__19_) );
INVX1 INVX1_966 ( .A(count_instr_20_), .Y(_1297_) );
NAND3X1 NAND3X1_75 ( .A(count_instr_16_), .B(count_instr_17_), .C(count_instr_18_), .Y(_1298_) );
NOR2X1 NOR2X1_1037 ( .A(_1294_), .B(_1298_), .Y(_1299_) );
NAND2X1 NAND2X1_762 ( .A(_1299_), .B(_1285_), .Y(_1300_) );
NOR2X1 NOR2X1_1038 ( .A(_10123__bF_buf0), .B(_1300_), .Y(_1301_) );
INVX1 INVX1_967 ( .A(_1301_), .Y(_1302_) );
NOR2X1 NOR2X1_1039 ( .A(_1297_), .B(_1302_), .Y(_1303_) );
OAI21X1 OAI21X1_2410 ( .A(_1301_), .B(count_instr_20_), .C(resetn_bF_buf1), .Y(_1304_) );
NOR2X1 NOR2X1_1040 ( .A(_1304_), .B(_1303_), .Y(_1__20_) );
INVX1 INVX1_968 ( .A(count_instr_21_), .Y(_1305_) );
INVX1 INVX1_969 ( .A(_1303_), .Y(_1306_) );
NOR2X1 NOR2X1_1041 ( .A(_1297_), .B(_1305_), .Y(_1307_) );
INVX1 INVX1_970 ( .A(_1307_), .Y(_1308_) );
OAI21X1 OAI21X1_2411 ( .A(_1302_), .B(_1308_), .C(resetn_bF_buf0), .Y(_1309_) );
AOI21X1 AOI21X1_824 ( .A(_1305_), .B(_1306_), .C(_1309_), .Y(_1__21_) );
NOR2X1 NOR2X1_1042 ( .A(_1308_), .B(_1302_), .Y(_1310_) );
OAI21X1 OAI21X1_2412 ( .A(_1310_), .B(count_instr_22_), .C(resetn_bF_buf11), .Y(_1311_) );
AOI21X1 AOI21X1_825 ( .A(count_instr_22_), .B(_1310_), .C(_1311_), .Y(_1__22_) );
AOI21X1 AOI21X1_826 ( .A(count_instr_22_), .B(_1310_), .C(count_instr_23_), .Y(_1312_) );
INVX1 INVX1_971 ( .A(_1310_), .Y(_1313_) );
NAND2X1 NAND2X1_763 ( .A(count_instr_22_), .B(count_instr_23_), .Y(_1314_) );
OAI21X1 OAI21X1_2413 ( .A(_1313_), .B(_1314_), .C(resetn_bF_buf10), .Y(_1315_) );
NOR2X1 NOR2X1_1043 ( .A(_1312_), .B(_1315_), .Y(_1__23_) );
OAI21X1 OAI21X1_2414 ( .A(_1313_), .B(_1314_), .C(count_instr_24_), .Y(_1316_) );
INVX1 INVX1_972 ( .A(count_instr_24_), .Y(_1317_) );
INVX1 INVX1_973 ( .A(_1314_), .Y(_1318_) );
NAND3X1 NAND3X1_76 ( .A(_1317_), .B(_1318_), .C(_1310_), .Y(_1319_) );
AOI21X1 AOI21X1_827 ( .A(_1319_), .B(_1316_), .C(_4426__bF_buf0), .Y(_1__24_) );
NAND2X1 NAND2X1_764 ( .A(_1318_), .B(_1307_), .Y(_1320_) );
NOR2X1 NOR2X1_1044 ( .A(_1320_), .B(_1300_), .Y(_1321_) );
INVX1 INVX1_974 ( .A(_1321_), .Y(_1322_) );
NAND2X1 NAND2X1_765 ( .A(count_instr_24_), .B(_10099__bF_buf1), .Y(_1323_) );
NOR2X1 NOR2X1_1045 ( .A(_1323_), .B(_1322_), .Y(_1324_) );
NOR2X1 NOR2X1_1046 ( .A(count_instr_25_), .B(_1324_), .Y(_1325_) );
AND2X2 AND2X2_186 ( .A(_1324_), .B(count_instr_25_), .Y(_1326_) );
NOR2X1 NOR2X1_1047 ( .A(_1325_), .B(_1326_), .Y(_1327_) );
AND2X2 AND2X2_187 ( .A(_1327_), .B(resetn_bF_buf9), .Y(_1__25_) );
XNOR2X1 XNOR2X1_47 ( .A(_1326_), .B(count_instr_26_), .Y(_1328_) );
NOR2X1 NOR2X1_1048 ( .A(_4426__bF_buf11), .B(_1328_), .Y(_1__26_) );
INVX1 INVX1_975 ( .A(count_instr_27_), .Y(_1329_) );
AND2X2 AND2X2_188 ( .A(count_instr_24_), .B(count_instr_25_), .Y(_1330_) );
NAND2X1 NAND2X1_766 ( .A(count_instr_26_), .B(_1330_), .Y(_1331_) );
NOR2X1 NOR2X1_1049 ( .A(_1331_), .B(_10123__bF_buf4), .Y(_1332_) );
AND2X2 AND2X2_189 ( .A(_1321_), .B(_1332_), .Y(_1333_) );
INVX1 INVX1_976 ( .A(_1333_), .Y(_1334_) );
OAI21X1 OAI21X1_2415 ( .A(_1334_), .B(_1329_), .C(resetn_bF_buf8), .Y(_1335_) );
AOI21X1 AOI21X1_828 ( .A(_1329_), .B(_1334_), .C(_1335_), .Y(_1__27_) );
NOR2X1 NOR2X1_1050 ( .A(_1329_), .B(_1331_), .Y(_1336_) );
NAND2X1 NAND2X1_767 ( .A(_1336_), .B(_1321_), .Y(_1337_) );
NOR2X1 NOR2X1_1051 ( .A(_10123__bF_buf3), .B(_1337_), .Y(_1338_) );
OAI21X1 OAI21X1_2416 ( .A(_1338_), .B(count_instr_28_), .C(resetn_bF_buf7), .Y(_1339_) );
AOI21X1 AOI21X1_829 ( .A(count_instr_28_), .B(_1338_), .C(_1339_), .Y(_1__28_) );
INVX1 INVX1_977 ( .A(count_instr_29_), .Y(_1340_) );
NAND2X1 NAND2X1_768 ( .A(count_instr_28_), .B(_1338_), .Y(_1341_) );
OAI21X1 OAI21X1_2417 ( .A(_1341_), .B(_1340_), .C(resetn_bF_buf6), .Y(_1342_) );
AOI21X1 AOI21X1_830 ( .A(_1340_), .B(_1341_), .C(_1342_), .Y(_1__29_) );
AND2X2 AND2X2_190 ( .A(count_instr_28_), .B(count_instr_29_), .Y(_1343_) );
NAND2X1 NAND2X1_769 ( .A(count_instr_30_), .B(_1343_), .Y(_1344_) );
INVX1 INVX1_978 ( .A(_1344_), .Y(_1345_) );
NOR2X1 NOR2X1_1052 ( .A(_1340_), .B(_1341_), .Y(_1346_) );
OAI21X1 OAI21X1_2418 ( .A(_1346_), .B(count_instr_30_), .C(resetn_bF_buf5), .Y(_1347_) );
AOI21X1 AOI21X1_831 ( .A(_1338_), .B(_1345_), .C(_1347_), .Y(_1__30_) );
AOI21X1 AOI21X1_832 ( .A(_1345_), .B(_1338_), .C(count_instr_31_), .Y(_1348_) );
INVX1 INVX1_979 ( .A(_1338_), .Y(_1349_) );
INVX1 INVX1_980 ( .A(count_instr_31_), .Y(_1350_) );
NOR2X1 NOR2X1_1053 ( .A(_1350_), .B(_1344_), .Y(_1351_) );
INVX1 INVX1_981 ( .A(_1351_), .Y(_1352_) );
OAI21X1 OAI21X1_2419 ( .A(_1349_), .B(_1352_), .C(resetn_bF_buf4), .Y(_1353_) );
NOR2X1 NOR2X1_1054 ( .A(_1348_), .B(_1353_), .Y(_1__31_) );
NOR2X1 NOR2X1_1055 ( .A(_1352_), .B(_1349_), .Y(_1354_) );
OAI21X1 OAI21X1_2420 ( .A(_1354_), .B(count_instr_32_), .C(resetn_bF_buf3), .Y(_1355_) );
AOI21X1 AOI21X1_833 ( .A(count_instr_32_), .B(_1354_), .C(_1355_), .Y(_1__32_) );
AOI21X1 AOI21X1_834 ( .A(count_instr_32_), .B(_1354_), .C(count_instr_33_), .Y(_1356_) );
NAND2X1 NAND2X1_770 ( .A(_1351_), .B(_1338_), .Y(_1357_) );
NAND2X1 NAND2X1_771 ( .A(count_instr_32_), .B(count_instr_33_), .Y(_1358_) );
OAI21X1 OAI21X1_2421 ( .A(_1357_), .B(_1358_), .C(resetn_bF_buf2), .Y(_1359_) );
NOR2X1 NOR2X1_1056 ( .A(_1359_), .B(_1356_), .Y(_1__33_) );
NOR2X1 NOR2X1_1057 ( .A(_1358_), .B(_1357_), .Y(_1360_) );
OAI21X1 OAI21X1_2422 ( .A(_1360_), .B(count_instr_34_), .C(resetn_bF_buf1), .Y(_1361_) );
AOI21X1 AOI21X1_835 ( .A(count_instr_34_), .B(_1360_), .C(_1361_), .Y(_1__34_) );
INVX1 INVX1_982 ( .A(count_instr_35_), .Y(_1362_) );
NAND2X1 NAND2X1_772 ( .A(count_instr_34_), .B(_1360_), .Y(_1363_) );
NAND2X1 NAND2X1_773 ( .A(count_instr_34_), .B(count_instr_35_), .Y(_1364_) );
NOR2X1 NOR2X1_1058 ( .A(_1358_), .B(_1364_), .Y(_1365_) );
INVX1 INVX1_983 ( .A(_1365_), .Y(_1366_) );
OAI21X1 OAI21X1_2423 ( .A(_1357_), .B(_1366_), .C(resetn_bF_buf0), .Y(_1367_) );
AOI21X1 AOI21X1_836 ( .A(_1362_), .B(_1363_), .C(_1367_), .Y(_1__35_) );
INVX1 INVX1_984 ( .A(count_instr_36_), .Y(_1368_) );
NOR2X1 NOR2X1_1059 ( .A(_1352_), .B(_1337_), .Y(_1369_) );
NAND3X1 NAND3X1_77 ( .A(_10099__bF_buf0), .B(_1365_), .C(_1369_), .Y(_1370_) );
OAI21X1 OAI21X1_2424 ( .A(_1370_), .B(_1368_), .C(resetn_bF_buf11), .Y(_1371_) );
AOI21X1 AOI21X1_837 ( .A(_1368_), .B(_1370_), .C(_1371_), .Y(_1__36_) );
INVX1 INVX1_985 ( .A(count_instr_37_), .Y(_1372_) );
NAND2X1 NAND2X1_774 ( .A(_1365_), .B(_1354_), .Y(_1373_) );
OR2X2 OR2X2_37 ( .A(_1373_), .B(_1368_), .Y(_1374_) );
NOR2X1 NOR2X1_1060 ( .A(_1368_), .B(_1372_), .Y(_1375_) );
INVX1 INVX1_986 ( .A(_1375_), .Y(_1376_) );
OAI21X1 OAI21X1_2425 ( .A(_1373_), .B(_1376_), .C(resetn_bF_buf10), .Y(_1377_) );
AOI21X1 AOI21X1_838 ( .A(_1372_), .B(_1374_), .C(_1377_), .Y(_1__37_) );
NOR2X1 NOR2X1_1061 ( .A(_1376_), .B(_1373_), .Y(_1378_) );
OAI21X1 OAI21X1_2426 ( .A(_1378_), .B(count_instr_38_), .C(resetn_bF_buf9), .Y(_1379_) );
AOI21X1 AOI21X1_839 ( .A(count_instr_38_), .B(_1378_), .C(_1379_), .Y(_1__38_) );
INVX1 INVX1_987 ( .A(count_instr_39_), .Y(_1380_) );
NAND2X1 NAND2X1_775 ( .A(count_instr_38_), .B(_1378_), .Y(_1381_) );
XNOR2X1 XNOR2X1_48 ( .A(_1381_), .B(_1380_), .Y(_1382_) );
NOR2X1 NOR2X1_1062 ( .A(_4426__bF_buf10), .B(_1382_), .Y(_1__39_) );
NAND2X1 NAND2X1_776 ( .A(count_instr_38_), .B(count_instr_39_), .Y(_1383_) );
NOR2X1 NOR2X1_1063 ( .A(_1383_), .B(_1376_), .Y(_1384_) );
NAND3X1 NAND3X1_78 ( .A(_1351_), .B(_1365_), .C(_1384_), .Y(_1385_) );
NOR2X1 NOR2X1_1064 ( .A(_1385_), .B(_1349_), .Y(_1386_) );
OAI21X1 OAI21X1_2427 ( .A(_1386_), .B(count_instr_40_), .C(resetn_bF_buf8), .Y(_1387_) );
AOI21X1 AOI21X1_840 ( .A(count_instr_40_), .B(_1386_), .C(_1387_), .Y(_1__40_) );
INVX1 INVX1_988 ( .A(count_instr_41_), .Y(_1388_) );
NAND3X1 NAND3X1_79 ( .A(_1365_), .B(_1384_), .C(_1369_), .Y(_1389_) );
NOR2X1 NOR2X1_1065 ( .A(_10123__bF_buf2), .B(_1389_), .Y(_1390_) );
AND2X2 AND2X2_191 ( .A(_1390_), .B(count_instr_40_), .Y(_1391_) );
INVX1 INVX1_989 ( .A(_1391_), .Y(_1392_) );
INVX1 INVX1_990 ( .A(count_instr_40_), .Y(_1393_) );
NOR2X1 NOR2X1_1066 ( .A(_1393_), .B(_1388_), .Y(_1394_) );
NAND2X1 NAND2X1_777 ( .A(_1394_), .B(_1386_), .Y(_1395_) );
NAND2X1 NAND2X1_778 ( .A(resetn_bF_buf7), .B(_1395_), .Y(_1396_) );
AOI21X1 AOI21X1_841 ( .A(_1388_), .B(_1392_), .C(_1396_), .Y(_1__41_) );
INVX1 INVX1_991 ( .A(count_instr_42_), .Y(_1397_) );
NOR2X1 NOR2X1_1067 ( .A(_1397_), .B(_1395_), .Y(_1398_) );
OAI21X1 OAI21X1_2428 ( .A(_1392_), .B(_1388_), .C(_1397_), .Y(_1399_) );
NAND2X1 NAND2X1_779 ( .A(resetn_bF_buf6), .B(_1399_), .Y(_1400_) );
NOR2X1 NOR2X1_1068 ( .A(_1398_), .B(_1400_), .Y(_1__42_) );
NOR2X1 NOR2X1_1069 ( .A(count_instr_43_), .B(_1398_), .Y(_1401_) );
INVX1 INVX1_992 ( .A(count_instr_43_), .Y(_1402_) );
NAND2X1 NAND2X1_780 ( .A(count_instr_42_), .B(_1394_), .Y(_1403_) );
NOR2X1 NOR2X1_1070 ( .A(_1402_), .B(_1403_), .Y(_1404_) );
NAND2X1 NAND2X1_781 ( .A(_1404_), .B(_1386_), .Y(_1405_) );
NAND2X1 NAND2X1_782 ( .A(resetn_bF_buf5), .B(_1405_), .Y(_1406_) );
NOR2X1 NOR2X1_1071 ( .A(_1406_), .B(_1401_), .Y(_1__43_) );
INVX1 INVX1_993 ( .A(count_instr_44_), .Y(_1407_) );
NOR2X1 NOR2X1_1072 ( .A(_1407_), .B(_1405_), .Y(_1408_) );
INVX1 INVX1_994 ( .A(_1405_), .Y(_1409_) );
OAI21X1 OAI21X1_2429 ( .A(_1409_), .B(count_instr_44_), .C(resetn_bF_buf4), .Y(_1410_) );
NOR2X1 NOR2X1_1073 ( .A(_1408_), .B(_1410_), .Y(_1__44_) );
OAI21X1 OAI21X1_2430 ( .A(_1405_), .B(_1407_), .C(count_instr_45_), .Y(_1411_) );
INVX1 INVX1_995 ( .A(count_instr_45_), .Y(_1412_) );
NAND2X1 NAND2X1_783 ( .A(_1412_), .B(_1408_), .Y(_1413_) );
AOI21X1 AOI21X1_842 ( .A(_1411_), .B(_1413_), .C(_4426__bF_buf9), .Y(_1__45_) );
INVX1 INVX1_996 ( .A(_1404_), .Y(_1414_) );
NOR2X1 NOR2X1_1074 ( .A(_1414_), .B(_1389_), .Y(_1415_) );
NOR2X1 NOR2X1_1075 ( .A(_1407_), .B(_1412_), .Y(_1416_) );
NAND2X1 NAND2X1_784 ( .A(_1416_), .B(_1415_), .Y(_1417_) );
NOR2X1 NOR2X1_1076 ( .A(_10123__bF_buf1), .B(_1417_), .Y(_1418_) );
NOR2X1 NOR2X1_1077 ( .A(count_instr_46_), .B(_1418_), .Y(_1419_) );
NAND2X1 NAND2X1_785 ( .A(count_instr_46_), .B(_1418_), .Y(_1420_) );
NAND2X1 NAND2X1_786 ( .A(resetn_bF_buf3), .B(_1420_), .Y(_1421_) );
NOR2X1 NOR2X1_1078 ( .A(_1419_), .B(_1421_), .Y(_1__46_) );
INVX1 INVX1_997 ( .A(count_instr_47_), .Y(_1422_) );
XNOR2X1 XNOR2X1_49 ( .A(_1420_), .B(_1422_), .Y(_1423_) );
NOR2X1 NOR2X1_1079 ( .A(_4426__bF_buf8), .B(_1423_), .Y(_1__47_) );
NOR2X1 NOR2X1_1080 ( .A(_1414_), .B(_1385_), .Y(_1424_) );
INVX1 INVX1_998 ( .A(count_instr_46_), .Y(_1425_) );
NOR2X1 NOR2X1_1081 ( .A(_1425_), .B(_1422_), .Y(_1426_) );
AND2X2 AND2X2_192 ( .A(_10099__bF_buf3), .B(_1426_), .Y(_1427_) );
NAND3X1 NAND3X1_80 ( .A(_1416_), .B(_1427_), .C(_1424_), .Y(_1428_) );
NOR2X1 NOR2X1_1082 ( .A(_1428_), .B(_1337_), .Y(_1429_) );
OAI21X1 OAI21X1_2431 ( .A(_1429_), .B(count_instr_48_), .C(resetn_bF_buf2), .Y(_1430_) );
AOI21X1 AOI21X1_843 ( .A(count_instr_48_), .B(_1429_), .C(_1430_), .Y(_1__48_) );
AOI21X1 AOI21X1_844 ( .A(count_instr_48_), .B(_1429_), .C(count_instr_49_), .Y(_1431_) );
INVX1 INVX1_999 ( .A(count_instr_48_), .Y(_1432_) );
INVX1 INVX1_1000 ( .A(count_instr_49_), .Y(_1433_) );
NOR2X1 NOR2X1_1083 ( .A(_1432_), .B(_1433_), .Y(_1434_) );
NAND2X1 NAND2X1_787 ( .A(_1434_), .B(_1429_), .Y(_1435_) );
NAND2X1 NAND2X1_788 ( .A(resetn_bF_buf1), .B(_1435_), .Y(_1436_) );
NOR2X1 NOR2X1_1084 ( .A(_1431_), .B(_1436_), .Y(_1__49_) );
INVX1 INVX1_1001 ( .A(count_instr_50_), .Y(_1437_) );
NAND3X1 NAND3X1_81 ( .A(_1416_), .B(_1426_), .C(_1415_), .Y(_1438_) );
NOR2X1 NOR2X1_1085 ( .A(_10123__bF_buf0), .B(_1438_), .Y(_1439_) );
NAND2X1 NAND2X1_789 ( .A(count_instr_50_), .B(_1434_), .Y(_1440_) );
INVX1 INVX1_1002 ( .A(_1440_), .Y(_1441_) );
NAND2X1 NAND2X1_790 ( .A(_1441_), .B(_1439_), .Y(_1442_) );
INVX1 INVX1_1003 ( .A(_1442_), .Y(_1443_) );
AOI21X1 AOI21X1_845 ( .A(_1437_), .B(_1435_), .C(_1443_), .Y(_1444_) );
AND2X2 AND2X2_193 ( .A(_1444_), .B(resetn_bF_buf0), .Y(_1__50_) );
INVX1 INVX1_1004 ( .A(count_instr_51_), .Y(_1445_) );
NOR2X1 NOR2X1_1086 ( .A(_1445_), .B(_1442_), .Y(_1446_) );
OAI21X1 OAI21X1_2432 ( .A(_1443_), .B(count_instr_51_), .C(resetn_bF_buf11), .Y(_1447_) );
NOR2X1 NOR2X1_1087 ( .A(_1446_), .B(_1447_), .Y(_1__51_) );
OAI21X1 OAI21X1_2433 ( .A(_1442_), .B(_1445_), .C(count_instr_52_), .Y(_1448_) );
INVX1 INVX1_1005 ( .A(count_instr_52_), .Y(_1449_) );
NAND2X1 NAND2X1_791 ( .A(_1449_), .B(_1446_), .Y(_1450_) );
AOI21X1 AOI21X1_846 ( .A(_1448_), .B(_1450_), .C(_4426__bF_buf7), .Y(_1__52_) );
INVX1 INVX1_1006 ( .A(count_instr_53_), .Y(_1451_) );
NOR2X1 NOR2X1_1088 ( .A(_1445_), .B(_1440_), .Y(_1452_) );
NAND2X1 NAND2X1_792 ( .A(count_instr_52_), .B(_1452_), .Y(_1453_) );
INVX1 INVX1_1007 ( .A(_1453_), .Y(_1454_) );
NAND2X1 NAND2X1_793 ( .A(_1454_), .B(_1439_), .Y(_1455_) );
OAI21X1 OAI21X1_2434 ( .A(_1455_), .B(_1451_), .C(resetn_bF_buf10), .Y(_1456_) );
AOI21X1 AOI21X1_847 ( .A(_1451_), .B(_1455_), .C(_1456_), .Y(_1__53_) );
NOR2X1 NOR2X1_1089 ( .A(_1451_), .B(_1455_), .Y(_1457_) );
NAND2X1 NAND2X1_794 ( .A(count_instr_54_), .B(_1457_), .Y(_1458_) );
INVX1 INVX1_1008 ( .A(_1458_), .Y(_1459_) );
OAI21X1 OAI21X1_2435 ( .A(_1457_), .B(count_instr_54_), .C(resetn_bF_buf9), .Y(_1460_) );
NOR2X1 NOR2X1_1090 ( .A(_1460_), .B(_1459_), .Y(_1__54_) );
INVX1 INVX1_1009 ( .A(count_instr_55_), .Y(_1461_) );
NOR2X1 NOR2X1_1091 ( .A(_1461_), .B(_1458_), .Y(_1462_) );
OAI21X1 OAI21X1_2436 ( .A(_1459_), .B(count_instr_55_), .C(resetn_bF_buf8), .Y(_1463_) );
NOR2X1 NOR2X1_1092 ( .A(_1462_), .B(_1463_), .Y(_1__55_) );
OAI21X1 OAI21X1_2437 ( .A(_1458_), .B(_1461_), .C(count_instr_56_), .Y(_1464_) );
INVX1 INVX1_1010 ( .A(count_instr_56_), .Y(_1465_) );
NAND2X1 NAND2X1_795 ( .A(_1465_), .B(_1462_), .Y(_1466_) );
AOI21X1 AOI21X1_848 ( .A(_1464_), .B(_1466_), .C(_4426__bF_buf6), .Y(_1__56_) );
NAND3X1 NAND3X1_82 ( .A(count_instr_53_), .B(count_instr_54_), .C(_1454_), .Y(_1467_) );
NOR2X1 NOR2X1_1093 ( .A(_1461_), .B(_1467_), .Y(_1468_) );
NAND2X1 NAND2X1_796 ( .A(count_instr_56_), .B(_1468_), .Y(_1469_) );
INVX1 INVX1_1011 ( .A(_1469_), .Y(_1470_) );
NAND2X1 NAND2X1_797 ( .A(_1429_), .B(_1470_), .Y(_1471_) );
INVX1 INVX1_1012 ( .A(_1471_), .Y(_1472_) );
AND2X2 AND2X2_194 ( .A(_1472_), .B(count_instr_57_), .Y(_1473_) );
OAI21X1 OAI21X1_2438 ( .A(_1472_), .B(count_instr_57_), .C(resetn_bF_buf7), .Y(_1474_) );
NOR2X1 NOR2X1_1094 ( .A(_1474_), .B(_1473_), .Y(_1__57_) );
AND2X2 AND2X2_195 ( .A(_1473_), .B(count_instr_58_), .Y(_1475_) );
OAI21X1 OAI21X1_2439 ( .A(_1473_), .B(count_instr_58_), .C(resetn_bF_buf6), .Y(_1476_) );
NOR2X1 NOR2X1_1095 ( .A(_1476_), .B(_1475_), .Y(_1__58_) );
AND2X2 AND2X2_196 ( .A(_1475_), .B(count_instr_59_), .Y(_1477_) );
OAI21X1 OAI21X1_2440 ( .A(_1475_), .B(count_instr_59_), .C(resetn_bF_buf5), .Y(_1478_) );
NOR2X1 NOR2X1_1096 ( .A(_1478_), .B(_1477_), .Y(_1__59_) );
INVX1 INVX1_1013 ( .A(count_instr_60_), .Y(_1479_) );
OR2X2 OR2X2_38 ( .A(_1477_), .B(_1479_), .Y(_1480_) );
NAND2X1 NAND2X1_798 ( .A(_1479_), .B(_1477_), .Y(_1481_) );
AOI21X1 AOI21X1_849 ( .A(_1481_), .B(_1480_), .C(_4426__bF_buf5), .Y(_1__60_) );
INVX1 INVX1_1014 ( .A(count_instr_61_), .Y(_1482_) );
NAND2X1 NAND2X1_799 ( .A(count_instr_57_), .B(count_instr_58_), .Y(_1483_) );
NAND2X1 NAND2X1_800 ( .A(count_instr_59_), .B(count_instr_60_), .Y(_1484_) );
NOR2X1 NOR2X1_1097 ( .A(_1483_), .B(_1484_), .Y(_1485_) );
NAND2X1 NAND2X1_801 ( .A(_1485_), .B(_1472_), .Y(_1486_) );
OAI21X1 OAI21X1_2441 ( .A(_1486_), .B(_1482_), .C(resetn_bF_buf4), .Y(_1487_) );
AOI21X1 AOI21X1_850 ( .A(_1482_), .B(_1486_), .C(_1487_), .Y(_1__61_) );
OAI21X1 OAI21X1_2442 ( .A(_1486_), .B(_1482_), .C(count_instr_62_), .Y(_1488_) );
INVX1 INVX1_1015 ( .A(count_instr_62_), .Y(_1489_) );
NOR2X1 NOR2X1_1098 ( .A(_1482_), .B(_1486_), .Y(_1490_) );
NAND2X1 NAND2X1_802 ( .A(_1489_), .B(_1490_), .Y(_1491_) );
AOI21X1 AOI21X1_851 ( .A(_1488_), .B(_1491_), .C(_4426__bF_buf4), .Y(_1__62_) );
NAND3X1 NAND3X1_83 ( .A(count_instr_61_), .B(count_instr_62_), .C(_1485_), .Y(_1492_) );
NOR2X1 NOR2X1_1099 ( .A(_1492_), .B(_1471_), .Y(_1493_) );
OAI21X1 OAI21X1_2443 ( .A(_1493_), .B(count_instr_63_), .C(resetn_bF_buf3), .Y(_1494_) );
AOI21X1 AOI21X1_852 ( .A(count_instr_63_), .B(_1493_), .C(_1494_), .Y(_1__63_) );
INVX1 INVX1_1016 ( .A(mem_rdata[19]), .Y(_1495_) );
NAND2X1 NAND2X1_803 ( .A(mem_rdata_q_19_), .B(_4439__bF_buf0), .Y(_1496_) );
OAI21X1 OAI21X1_2444 ( .A(_1495_), .B(_4439__bF_buf6), .C(_1496_), .Y(mem_rdata_latched_19_) );
NAND2X1 NAND2X1_804 ( .A(mem_rdata_latched_19_), .B(_4985__bF_buf7), .Y(_1497_) );
OAI21X1 OAI21X1_2445 ( .A(_7552__bF_buf5), .B(_4985__bF_buf6), .C(_1497_), .Y(_5__4_) );
INVX1 INVX1_1017 ( .A(mem_rdata[30]), .Y(_1498_) );
NAND2X1 NAND2X1_805 ( .A(mem_rdata_q_30_), .B(_4439__bF_buf5), .Y(_1499_) );
OAI21X1 OAI21X1_2446 ( .A(_1498_), .B(_4439__bF_buf4), .C(_1499_), .Y(mem_rdata_latched_30_) );
NAND2X1 NAND2X1_806 ( .A(mem_rdata_latched_30_), .B(_4985__bF_buf5), .Y(_1500_) );
OAI21X1 OAI21X1_2447 ( .A(_10288_), .B(_4985__bF_buf4), .C(_1500_), .Y(_3__10_) );
INVX1 INVX1_1018 ( .A(mem_rdata[27]), .Y(_1501_) );
NAND2X1 NAND2X1_807 ( .A(mem_rdata_q_27_), .B(_4439__bF_buf3), .Y(_1502_) );
OAI21X1 OAI21X1_2448 ( .A(_1501_), .B(_4439__bF_buf2), .C(_1502_), .Y(mem_rdata_latched_27_) );
NAND2X1 NAND2X1_808 ( .A(mem_rdata_latched_27_), .B(_4985__bF_buf3), .Y(_1503_) );
OAI21X1 OAI21X1_2449 ( .A(_10225_), .B(_4985__bF_buf2), .C(_1503_), .Y(_3__7_) );
INVX1 INVX1_1019 ( .A(mem_rdata[26]), .Y(_1504_) );
NAND2X1 NAND2X1_809 ( .A(mem_rdata_q_26_), .B(_4439__bF_buf1), .Y(_1505_) );
OAI21X1 OAI21X1_2450 ( .A(_1504_), .B(_4439__bF_buf0), .C(_1505_), .Y(mem_rdata_latched_26_) );
NAND2X1 NAND2X1_810 ( .A(mem_rdata_latched_26_), .B(_4985__bF_buf1), .Y(_1506_) );
OAI21X1 OAI21X1_2451 ( .A(_10213_), .B(_4985__bF_buf0), .C(_1506_), .Y(_3__6_) );
INVX1 INVX1_1020 ( .A(mem_rdata_q_21_), .Y(_1507_) );
NAND2X1 NAND2X1_811 ( .A(mem_rdata[21]), .B(_4542_), .Y(_1508_) );
OAI21X1 OAI21X1_2452 ( .A(_1507_), .B(_4542_), .C(_1508_), .Y(mem_rdata_latched_21_) );
NAND2X1 NAND2X1_812 ( .A(mem_rdata_latched_21_), .B(_4985__bF_buf8), .Y(_1509_) );
OAI21X1 OAI21X1_2453 ( .A(_10112_), .B(_4985__bF_buf7), .C(_1509_), .Y(_3__1_) );
INVX1 INVX1_1021 ( .A(mem_rdata_q_22_), .Y(_1510_) );
NAND2X1 NAND2X1_813 ( .A(mem_rdata[22]), .B(_4542_), .Y(_1511_) );
OAI21X1 OAI21X1_2454 ( .A(_1510_), .B(_4542_), .C(_1511_), .Y(mem_rdata_latched_22_) );
NAND2X1 NAND2X1_814 ( .A(mem_rdata_latched_22_), .B(_4985__bF_buf6), .Y(_1512_) );
OAI21X1 OAI21X1_2455 ( .A(_10133_), .B(_4985__bF_buf5), .C(_1512_), .Y(_3__2_) );
INVX1 INVX1_1022 ( .A(mem_rdata[23]), .Y(_1513_) );
NAND2X1 NAND2X1_815 ( .A(mem_rdata_q_23_), .B(_4439__bF_buf6), .Y(_1514_) );
OAI21X1 OAI21X1_2456 ( .A(_1513_), .B(_4439__bF_buf5), .C(_1514_), .Y(mem_rdata_latched_23_) );
NAND2X1 NAND2X1_816 ( .A(mem_rdata_latched_23_), .B(_4985__bF_buf4), .Y(_1515_) );
OAI21X1 OAI21X1_2457 ( .A(_10150_), .B(_4985__bF_buf3), .C(_1515_), .Y(_3__3_) );
INVX1 INVX1_1023 ( .A(mem_rdata[25]), .Y(_1516_) );
NAND2X1 NAND2X1_817 ( .A(mem_rdata_q_25_), .B(_4439__bF_buf4), .Y(_1517_) );
OAI21X1 OAI21X1_2458 ( .A(_1516_), .B(_4439__bF_buf3), .C(_1517_), .Y(mem_rdata_latched_25_) );
NAND2X1 NAND2X1_818 ( .A(mem_rdata_latched_25_), .B(_4985__bF_buf2), .Y(_1518_) );
OAI21X1 OAI21X1_2459 ( .A(_10190_), .B(_4985__bF_buf1), .C(_1518_), .Y(_3__5_) );
INVX1 INVX1_1024 ( .A(mem_rdata[28]), .Y(_1519_) );
NAND2X1 NAND2X1_819 ( .A(mem_rdata_q_28_), .B(_4439__bF_buf2), .Y(_1520_) );
OAI21X1 OAI21X1_2460 ( .A(_1519_), .B(_4439__bF_buf1), .C(_1520_), .Y(mem_rdata_latched_28_) );
NAND2X1 NAND2X1_820 ( .A(mem_rdata_latched_28_), .B(_4985__bF_buf0), .Y(_1521_) );
OAI21X1 OAI21X1_2461 ( .A(_10339_), .B(_4985__bF_buf8), .C(_1521_), .Y(_3__8_) );
INVX1 INVX1_1025 ( .A(mem_rdata[29]), .Y(_1522_) );
NAND2X1 NAND2X1_821 ( .A(mem_rdata_q_29_), .B(_4439__bF_buf0), .Y(_1523_) );
OAI21X1 OAI21X1_2462 ( .A(_1522_), .B(_4439__bF_buf6), .C(_1523_), .Y(mem_rdata_latched_29_) );
NAND2X1 NAND2X1_822 ( .A(mem_rdata_latched_29_), .B(_4985__bF_buf7), .Y(_1524_) );
OAI21X1 OAI21X1_2463 ( .A(_10269_), .B(_4985__bF_buf6), .C(_1524_), .Y(_3__9_) );
INVX1 INVX1_1026 ( .A(mem_rdata[31]), .Y(_1525_) );
NAND2X1 NAND2X1_823 ( .A(mem_rdata_q_31_), .B(_4439__bF_buf5), .Y(_1526_) );
OAI21X1 OAI21X1_2464 ( .A(_1525_), .B(_4439__bF_buf4), .C(_1526_), .Y(mem_rdata_latched_31_) );
NAND2X1 NAND2X1_824 ( .A(mem_rdata_latched_31_), .B(_4985__bF_buf5), .Y(_1527_) );
OAI21X1 OAI21X1_2465 ( .A(_10519_), .B(_4985__bF_buf4), .C(_1527_), .Y(_3__20_) );
OAI21X1 OAI21X1_2466 ( .A(_10537_), .B(_4985__bF_buf3), .C(_1527_), .Y(_3__21_) );
OAI21X1 OAI21X1_2467 ( .A(_10559_), .B(_4985__bF_buf2), .C(_1527_), .Y(_3__22_) );
OAI21X1 OAI21X1_2468 ( .A(_10579_), .B(_4985__bF_buf1), .C(_1527_), .Y(_3__23_) );
OAI21X1 OAI21X1_2469 ( .A(_10612_), .B(_4985__bF_buf0), .C(_1527_), .Y(_3__24_) );
OAI21X1 OAI21X1_2470 ( .A(_10632_), .B(_4985__bF_buf8), .C(_1527_), .Y(_3__25_) );
OAI21X1 OAI21X1_2471 ( .A(_10652_), .B(_4985__bF_buf7), .C(_1527_), .Y(_3__26_) );
OAI21X1 OAI21X1_2472 ( .A(_10670_), .B(_4985__bF_buf6), .C(_1527_), .Y(_3__27_) );
OAI21X1 OAI21X1_2473 ( .A(_10700_), .B(_4985__bF_buf5), .C(_1527_), .Y(_3__28_) );
OAI21X1 OAI21X1_2474 ( .A(_10716_), .B(_4985__bF_buf4), .C(_1527_), .Y(_3__29_) );
INVX1 INVX1_1027 ( .A(decoded_imm_uj_30_), .Y(_1528_) );
OAI21X1 OAI21X1_2475 ( .A(_1528_), .B(_4985__bF_buf3), .C(_1527_), .Y(_3__30_) );
OAI21X1 OAI21X1_2476 ( .A(_1169_), .B(_4985__bF_buf2), .C(_1527_), .Y(_3__31_) );
INVX1 INVX1_1028 ( .A(mem_rdata[24]), .Y(_1529_) );
NAND2X1 NAND2X1_825 ( .A(mem_rdata_q_24_), .B(_4439__bF_buf3), .Y(_1530_) );
OAI21X1 OAI21X1_2477 ( .A(_1529_), .B(_4439__bF_buf2), .C(_1530_), .Y(mem_rdata_latched_24_) );
NAND2X1 NAND2X1_826 ( .A(mem_rdata_latched_24_), .B(_4985__bF_buf1), .Y(_1531_) );
OAI21X1 OAI21X1_2478 ( .A(_10163_), .B(_4985__bF_buf0), .C(_1531_), .Y(_3__4_) );
INVX1 INVX1_1029 ( .A(mem_rdata[20]), .Y(_1532_) );
NAND2X1 NAND2X1_827 ( .A(mem_rdata_q_20_), .B(_4439__bF_buf1), .Y(_1533_) );
OAI21X1 OAI21X1_2479 ( .A(_1532_), .B(_4439__bF_buf0), .C(_1533_), .Y(mem_rdata_latched_20_) );
NAND2X1 NAND2X1_828 ( .A(mem_rdata_latched_20_), .B(_4985__bF_buf8), .Y(_1534_) );
OAI21X1 OAI21X1_2480 ( .A(_10313_), .B(_4985__bF_buf7), .C(_1534_), .Y(_3__11_) );
NOR2X1 NOR2X1_1100 ( .A(_10100_), .B(_4985__bF_buf6), .Y(_3__0_) );
INVX1 INVX1_1030 ( .A(mem_rdata[15]), .Y(_1535_) );
NAND2X1 NAND2X1_829 ( .A(mem_rdata_q_15_), .B(_4439__bF_buf6), .Y(_1536_) );
OAI21X1 OAI21X1_2481 ( .A(_1535_), .B(_4439__bF_buf5), .C(_1536_), .Y(mem_rdata_latched_15_) );
NAND2X1 NAND2X1_830 ( .A(mem_rdata_latched_15_), .B(_4985__bF_buf5), .Y(_1537_) );
OAI21X1 OAI21X1_2482 ( .A(_7569__bF_buf43), .B(_4985__bF_buf4), .C(_1537_), .Y(_5__0_) );
INVX1 INVX1_1031 ( .A(mem_rdata_q_16_), .Y(_1538_) );
NAND2X1 NAND2X1_831 ( .A(mem_rdata[16]), .B(_4542_), .Y(_1539_) );
OAI21X1 OAI21X1_2483 ( .A(_1538_), .B(_4542_), .C(_1539_), .Y(mem_rdata_latched_16_) );
NAND2X1 NAND2X1_832 ( .A(mem_rdata_latched_16_), .B(_4985__bF_buf3), .Y(_1540_) );
OAI21X1 OAI21X1_2484 ( .A(_7556__bF_buf17), .B(_4985__bF_buf2), .C(_1540_), .Y(_5__1_) );
INVX1 INVX1_1032 ( .A(mem_rdata[17]), .Y(_1541_) );
NAND2X1 NAND2X1_833 ( .A(mem_rdata_q_17_), .B(_4439__bF_buf4), .Y(_1542_) );
OAI21X1 OAI21X1_2485 ( .A(_1541_), .B(_4439__bF_buf3), .C(_1542_), .Y(mem_rdata_latched_17_) );
NAND2X1 NAND2X1_834 ( .A(mem_rdata_latched_17_), .B(_4985__bF_buf1), .Y(_1543_) );
OAI21X1 OAI21X1_2486 ( .A(_7560__bF_buf0), .B(_4985__bF_buf0), .C(_1543_), .Y(_5__2_) );
INVX1 INVX1_1033 ( .A(mem_rdata[18]), .Y(_1544_) );
NAND2X1 NAND2X1_835 ( .A(mem_rdata_q_18_), .B(_4439__bF_buf2), .Y(_1545_) );
OAI21X1 OAI21X1_2487 ( .A(_1544_), .B(_4439__bF_buf1), .C(_1545_), .Y(mem_rdata_latched_18_) );
NAND2X1 NAND2X1_836 ( .A(mem_rdata_latched_18_), .B(_4985__bF_buf8), .Y(_1546_) );
OAI21X1 OAI21X1_2488 ( .A(_7561__bF_buf3), .B(_4985__bF_buf7), .C(_1546_), .Y(_5__3_) );
NOR2X1 NOR2X1_1101 ( .A(decoder_pseudo_trigger_bF_buf3), .B(_4605__bF_buf5), .Y(_1547_) );
NOR2X1 NOR2X1_1102 ( .A(_57_), .B(_4510_), .Y(_1548_) );
NOR2X1 NOR2X1_1103 ( .A(_1547__bF_buf5), .B(_1548_), .Y(_58_) );
INVX1 INVX1_1034 ( .A(mem_rdata[0]), .Y(_1549_) );
NAND2X1 NAND2X1_837 ( .A(mem_rdata_q_0_), .B(_4439__bF_buf0), .Y(_1550_) );
OAI21X1 OAI21X1_2489 ( .A(_1549_), .B(_4439__bF_buf6), .C(_1550_), .Y(mem_rdata_latched_0_) );
INVX1 INVX1_1035 ( .A(mem_rdata[1]), .Y(_1551_) );
NAND2X1 NAND2X1_838 ( .A(mem_rdata_q_1_), .B(_4439__bF_buf5), .Y(_1552_) );
OAI21X1 OAI21X1_2490 ( .A(_1551_), .B(_4439__bF_buf4), .C(_1552_), .Y(mem_rdata_latched_1_) );
INVX1 INVX1_1036 ( .A(is_alu_reg_reg), .Y(_1553_) );
INVX1 INVX1_1037 ( .A(mem_rdata_latched_5_), .Y(_1554_) );
NAND2X1 NAND2X1_839 ( .A(_4548_), .B(mem_rdata_latched_4_), .Y(_1555_) );
NOR2X1 NOR2X1_1104 ( .A(_1555_), .B(_1554_), .Y(_1556_) );
NAND2X1 NAND2X1_840 ( .A(mem_rdata_latched_0_), .B(mem_rdata_latched_1_), .Y(_1557_) );
INVX1 INVX1_1038 ( .A(_1557_), .Y(_1558_) );
NOR2X1 NOR2X1_1105 ( .A(mem_rdata_latched_2_), .B(mem_rdata_latched_3_), .Y(_1559_) );
NAND2X1 NAND2X1_841 ( .A(_1558_), .B(_1559_), .Y(_1560_) );
INVX1 INVX1_1039 ( .A(_1560_), .Y(_1561_) );
NAND3X1 NAND3X1_84 ( .A(_1556_), .B(_1561_), .C(_4985__bF_buf6), .Y(_1562_) );
OAI21X1 OAI21X1_2491 ( .A(_1553_), .B(_4985__bF_buf5), .C(_1562_), .Y(_51_) );
INVX1 INVX1_1040 ( .A(is_alu_reg_imm), .Y(_1563_) );
NOR2X1 NOR2X1_1106 ( .A(mem_rdata_latched_5_), .B(_1555_), .Y(_1564_) );
NAND3X1 NAND3X1_85 ( .A(_1564_), .B(_1561_), .C(_4985__bF_buf4), .Y(_1565_) );
OAI21X1 OAI21X1_2492 ( .A(_1563_), .B(_4985__bF_buf3), .C(_1565_), .Y(_50_) );
INVX1 INVX1_1041 ( .A(_1547__bF_buf4), .Y(_1566_) );
NOR2X1 NOR2X1_1107 ( .A(_1553_), .B(_1566__bF_buf3), .Y(_1567_) );
INVX1 INVX1_1042 ( .A(_1567_), .Y(_1568_) );
NOR2X1 NOR2X1_1108 ( .A(mem_rdata_q_27_), .B(mem_rdata_q_26_), .Y(_1569_) );
INVX1 INVX1_1043 ( .A(_1569_), .Y(_1570_) );
NOR2X1 NOR2X1_1109 ( .A(mem_rdata_q_25_), .B(mem_rdata_q_28_), .Y(_1571_) );
NOR2X1 NOR2X1_1110 ( .A(mem_rdata_q_29_), .B(mem_rdata_q_31_), .Y(_1572_) );
NAND2X1 NAND2X1_842 ( .A(_1571_), .B(_1572_), .Y(_1573_) );
NOR2X1 NOR2X1_1111 ( .A(_1570_), .B(_1573_), .Y(_1574_) );
INVX1 INVX1_1044 ( .A(mem_rdata_q_14_), .Y(_1575_) );
INVX1 INVX1_1045 ( .A(mem_rdata_q_12_), .Y(_1576_) );
NOR2X1 NOR2X1_1112 ( .A(mem_rdata_q_13_), .B(_1576_), .Y(_1577_) );
INVX1 INVX1_1046 ( .A(_1577_), .Y(_1578_) );
AOI21X1 AOI21X1_853 ( .A(_1575_), .B(mem_rdata_q_30_), .C(_1578_), .Y(_1579_) );
NAND2X1 NAND2X1_843 ( .A(_1574_), .B(_1579_), .Y(_1580_) );
OAI22X1 OAI22X1_227 ( .A(_4572_), .B(_1547__bF_buf3), .C(_1580_), .D(_1568_), .Y(_60_) );
NOR2X1 NOR2X1_1113 ( .A(mem_rdata_latched_4_), .B(_1554_), .Y(_1581_) );
NOR2X1 NOR2X1_1114 ( .A(mem_rdata_latched_6_), .B(_1560_), .Y(_1582_) );
NAND3X1 NAND3X1_86 ( .A(_4985__bF_buf2), .B(_1581_), .C(_1582_), .Y(_1583_) );
OAI21X1 OAI21X1_2493 ( .A(_4592_), .B(_4985__bF_buf1), .C(_1583_), .Y(_59_) );
NOR2X1 NOR2X1_1115 ( .A(_1563_), .B(_1566__bF_buf2), .Y(_1584_) );
INVX1 INVX1_1047 ( .A(_1584_), .Y(_1585_) );
MUX2X1 MUX2X1_232 ( .A(instr_jalr), .B(is_jalr_addi_slti_sltiu_xori_ori_andi), .S(_1547__bF_buf2), .Y(_1586_) );
OAI21X1 OAI21X1_2494 ( .A(_1585_), .B(_1577_), .C(_1586_), .Y(_54_) );
OAI22X1 OAI22X1_228 ( .A(_4564_), .B(_1547__bF_buf1), .C(_1580_), .D(_1585_), .Y(_61_) );
INVX1 INVX1_1048 ( .A(_4985__bF_buf0), .Y(_1587_) );
NOR2X1 NOR2X1_1116 ( .A(mem_rdata_latched_4_), .B(mem_rdata_latched_5_), .Y(_1588_) );
NAND2X1 NAND2X1_844 ( .A(_1588_), .B(_1582_), .Y(_1589_) );
OAI21X1 OAI21X1_2495 ( .A(_4588_), .B(_4984_), .C(is_lb_lh_lw_lbu_lhu), .Y(_1590_) );
OAI21X1 OAI21X1_2496 ( .A(_1589_), .B(_1587_), .C(_1590_), .Y(_55_) );
NAND2X1 NAND2X1_845 ( .A(_5847_), .B(_1563_), .Y(_1591_) );
NOR2X1 NOR2X1_1117 ( .A(is_lb_lh_lw_lbu_lhu), .B(_1591_), .Y(_1592_) );
INVX1 INVX1_1049 ( .A(_1592_), .Y(_1593_) );
INVX1 INVX1_1050 ( .A(mem_rdata_q_7_), .Y(_1594_) );
INVX1 INVX1_1051 ( .A(_10101_), .Y(_1595_) );
OAI21X1 OAI21X1_2497 ( .A(_4592_), .B(_1594_), .C(_1595_), .Y(_1596_) );
AOI21X1 AOI21X1_854 ( .A(mem_rdata_q_20_), .B(_1593_), .C(_1596_), .Y(_1597_) );
OAI21X1 OAI21X1_2498 ( .A(_4605__bF_buf4), .B(decoder_pseudo_trigger_bF_buf2), .C(decoded_imm_0_), .Y(_1598_) );
OAI21X1 OAI21X1_2499 ( .A(_1597_), .B(_1566__bF_buf1), .C(_1598_), .Y(_2__0_) );
NOR2X1 NOR2X1_1118 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .Y(_1599_) );
NAND2X1 NAND2X1_846 ( .A(_1599_), .B(_1592_), .Y(_1600_) );
OAI21X1 OAI21X1_2500 ( .A(_1600_), .B(_57_), .C(_1547__bF_buf0), .Y(_1601_) );
OAI21X1 OAI21X1_2501 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(mem_rdata_q_8_), .Y(_1602_) );
OAI21X1 OAI21X1_2502 ( .A(_4499__bF_buf5), .B(_10112_), .C(_1602_), .Y(_1603_) );
AOI21X1 AOI21X1_855 ( .A(mem_rdata_q_21_), .B(_1593_), .C(_1603_), .Y(_1604_) );
OAI22X1 OAI22X1_229 ( .A(_7762_), .B(_1547__bF_buf5), .C(_1601__bF_buf4), .D(_1604_), .Y(_2__1_) );
OAI21X1 OAI21X1_2503 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(mem_rdata_q_9_), .Y(_1605_) );
OAI21X1 OAI21X1_2504 ( .A(_4499__bF_buf4), .B(_10133_), .C(_1605_), .Y(_1606_) );
AOI21X1 AOI21X1_856 ( .A(mem_rdata_q_22_), .B(_1593_), .C(_1606_), .Y(_1607_) );
OAI22X1 OAI22X1_230 ( .A(_7766_), .B(_1547__bF_buf4), .C(_1601__bF_buf3), .D(_1607_), .Y(_2__2_) );
OAI21X1 OAI21X1_2505 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(mem_rdata_q_10_), .Y(_1608_) );
OAI21X1 OAI21X1_2506 ( .A(_4499__bF_buf3), .B(_10150_), .C(_1608_), .Y(_1609_) );
AOI21X1 AOI21X1_857 ( .A(mem_rdata_q_23_), .B(_1593_), .C(_1609_), .Y(_1610_) );
OAI22X1 OAI22X1_231 ( .A(_7850_), .B(_1547__bF_buf3), .C(_1601__bF_buf2), .D(_1610_), .Y(_2__3_) );
OAI21X1 OAI21X1_2507 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(mem_rdata_q_11_), .Y(_1611_) );
OAI21X1 OAI21X1_2508 ( .A(_4499__bF_buf2), .B(_10163_), .C(_1611_), .Y(_1612_) );
AOI21X1 AOI21X1_858 ( .A(mem_rdata_q_24_), .B(_1593_), .C(_1612_), .Y(_1613_) );
OAI22X1 OAI22X1_232 ( .A(_7914_), .B(_1547__bF_buf2), .C(_1601__bF_buf1), .D(_1613_), .Y(_2__4_) );
AOI22X1 AOI22X1_106 ( .A(instr_jal_bF_buf1), .B(decoded_imm_uj_5_), .C(_1600_), .D(mem_rdata_q_25_), .Y(_1614_) );
OAI22X1 OAI22X1_233 ( .A(_7926_), .B(_1547__bF_buf1), .C(_1614_), .D(_1601__bF_buf0), .Y(_2__5_) );
AOI22X1 AOI22X1_107 ( .A(instr_jal_bF_buf0), .B(decoded_imm_uj_6_), .C(_1600_), .D(mem_rdata_q_26_), .Y(_1615_) );
OAI22X1 OAI22X1_234 ( .A(_8005_), .B(_1547__bF_buf0), .C(_1615_), .D(_1601__bF_buf4), .Y(_2__6_) );
AOI22X1 AOI22X1_108 ( .A(instr_jal_bF_buf6), .B(decoded_imm_uj_7_), .C(_1600_), .D(mem_rdata_q_27_), .Y(_1616_) );
OAI22X1 OAI22X1_235 ( .A(_8070_), .B(_1547__bF_buf5), .C(_1616_), .D(_1601__bF_buf3), .Y(_2__7_) );
AOI22X1 AOI22X1_109 ( .A(instr_jal_bF_buf5), .B(decoded_imm_uj_8_), .C(_1600_), .D(mem_rdata_q_28_), .Y(_1617_) );
OAI22X1 OAI22X1_236 ( .A(_8230_), .B(_1547__bF_buf4), .C(_1617_), .D(_1601__bF_buf2), .Y(_2__8_) );
AOI22X1 AOI22X1_110 ( .A(instr_jal_bF_buf4), .B(decoded_imm_uj_9_), .C(_1600_), .D(mem_rdata_q_29_), .Y(_1618_) );
OAI22X1 OAI22X1_237 ( .A(_8225_), .B(_1547__bF_buf3), .C(_1618_), .D(_1601__bF_buf1), .Y(_2__9_) );
AOI22X1 AOI22X1_111 ( .A(instr_jal_bF_buf3), .B(decoded_imm_uj_10_), .C(_1600_), .D(mem_rdata_q_30_), .Y(_1619_) );
OAI22X1 OAI22X1_238 ( .A(_8304_), .B(_1547__bF_buf2), .C(_1619_), .D(_1601__bF_buf0), .Y(_2__10_) );
OAI21X1 OAI21X1_2509 ( .A(_1591_), .B(is_lb_lh_lw_lbu_lhu), .C(mem_rdata_q_31_), .Y(_1620_) );
NAND2X1 NAND2X1_847 ( .A(is_sb_sh_sw), .B(mem_rdata_q_31_), .Y(_1621_) );
OAI21X1 OAI21X1_2510 ( .A(_4556_), .B(_1594_), .C(_1621_), .Y(_1622_) );
AOI21X1 AOI21X1_859 ( .A(instr_jal_bF_buf2), .B(decoded_imm_uj_11_), .C(_1622_), .Y(_1623_) );
AND2X2 AND2X2_197 ( .A(_1623_), .B(_1620_), .Y(_1624_) );
OAI22X1 OAI22X1_239 ( .A(_8459_), .B(_1547__bF_buf1), .C(_1601__bF_buf4), .D(_1624_), .Y(_2__11_) );
OAI21X1 OAI21X1_2511 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_12_), .Y(_1625_) );
OAI21X1 OAI21X1_2512 ( .A(is_sb_sh_sw), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(mem_rdata_q_31_), .Y(_1626_) );
AND2X2 AND2X2_198 ( .A(_1625_), .B(_1626_), .Y(_1627_) );
OAI21X1 OAI21X1_2513 ( .A(_4499__bF_buf1), .B(_10347_), .C(_1627_), .Y(_1628_) );
AOI21X1 AOI21X1_860 ( .A(mem_rdata_q_31_), .B(_1593_), .C(_1628_), .Y(_1629_) );
OAI22X1 OAI22X1_240 ( .A(_8465_), .B(_1547__bF_buf0), .C(_1601__bF_buf3), .D(_1629_), .Y(_2__12_) );
NAND2X1 NAND2X1_848 ( .A(_1626_), .B(_1620_), .Y(_1630_) );
INVX1 INVX1_1052 ( .A(mem_rdata_q_13_), .Y(_1631_) );
OAI22X1 OAI22X1_241 ( .A(_4499__bF_buf0), .B(_10360_), .C(_4500_), .D(_1631_), .Y(_1632_) );
NOR2X1 NOR2X1_1119 ( .A(_1632_), .B(_1630__bF_buf3), .Y(_1633_) );
OAI22X1 OAI22X1_242 ( .A(_8543_), .B(_1547__bF_buf5), .C(_1601__bF_buf2), .D(_1633_), .Y(_2__13_) );
OAI22X1 OAI22X1_243 ( .A(_4499__bF_buf5), .B(_10382_), .C(_4500_), .D(_1575_), .Y(_1634_) );
NOR2X1 NOR2X1_1120 ( .A(_1634_), .B(_1630__bF_buf2), .Y(_1635_) );
OAI22X1 OAI22X1_244 ( .A(_8623_), .B(_1547__bF_buf4), .C(_1601__bF_buf1), .D(_1635_), .Y(_2__14_) );
INVX1 INVX1_1053 ( .A(mem_rdata_q_15_), .Y(_1636_) );
OAI22X1 OAI22X1_245 ( .A(_4499__bF_buf4), .B(_10397_), .C(_4500_), .D(_1636_), .Y(_1637_) );
NOR2X1 NOR2X1_1121 ( .A(_1637_), .B(_1630__bF_buf1), .Y(_1638_) );
OAI22X1 OAI22X1_246 ( .A(_8775_), .B(_1547__bF_buf3), .C(_1601__bF_buf0), .D(_1638_), .Y(_2__15_) );
OAI22X1 OAI22X1_247 ( .A(_4499__bF_buf3), .B(_10433_), .C(_4500_), .D(_1538_), .Y(_1639_) );
NOR2X1 NOR2X1_1122 ( .A(_1639_), .B(_1630__bF_buf0), .Y(_1640_) );
OAI22X1 OAI22X1_248 ( .A(_8782_), .B(_1547__bF_buf2), .C(_1601__bF_buf4), .D(_1640_), .Y(_2__16_) );
OAI21X1 OAI21X1_2514 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_17_), .Y(_1641_) );
OAI21X1 OAI21X1_2515 ( .A(_4499__bF_buf2), .B(_10454_), .C(_1641_), .Y(_1642_) );
NOR2X1 NOR2X1_1123 ( .A(_1642_), .B(_1630__bF_buf3), .Y(_1643_) );
OAI22X1 OAI22X1_249 ( .A(_8868_), .B(_1547__bF_buf1), .C(_1601__bF_buf3), .D(_1643_), .Y(_2__17_) );
OAI21X1 OAI21X1_2516 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_18_), .Y(_1644_) );
OAI21X1 OAI21X1_2517 ( .A(_4499__bF_buf1), .B(_10470_), .C(_1644_), .Y(_1645_) );
NOR2X1 NOR2X1_1124 ( .A(_1645_), .B(_1630__bF_buf2), .Y(_1646_) );
OAI22X1 OAI22X1_250 ( .A(_8947_), .B(_1547__bF_buf0), .C(_1601__bF_buf2), .D(_1646_), .Y(_2__18_) );
INVX1 INVX1_1054 ( .A(decoded_imm_19_), .Y(_1647_) );
OAI21X1 OAI21X1_2518 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_19_), .Y(_1648_) );
OAI21X1 OAI21X1_2519 ( .A(_4499__bF_buf0), .B(_10490_), .C(_1648_), .Y(_1649_) );
NOR2X1 NOR2X1_1125 ( .A(_1649_), .B(_1630__bF_buf1), .Y(_1650_) );
OAI22X1 OAI22X1_251 ( .A(_1647_), .B(_1547__bF_buf5), .C(_1601__bF_buf1), .D(_1650_), .Y(_2__19_) );
OAI21X1 OAI21X1_2520 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_20_), .Y(_1651_) );
OAI21X1 OAI21X1_2521 ( .A(_4499__bF_buf5), .B(_10519_), .C(_1651_), .Y(_1652_) );
NOR2X1 NOR2X1_1126 ( .A(_1652_), .B(_1630__bF_buf0), .Y(_1653_) );
OAI22X1 OAI22X1_252 ( .A(_9107_), .B(_1547__bF_buf4), .C(_1601__bF_buf0), .D(_1653_), .Y(_2__20_) );
INVX1 INVX1_1055 ( .A(decoded_imm_21_), .Y(_1654_) );
OAI22X1 OAI22X1_253 ( .A(_4499__bF_buf4), .B(_10537_), .C(_4500_), .D(_1507_), .Y(_1655_) );
NOR2X1 NOR2X1_1127 ( .A(_1655_), .B(_1630__bF_buf3), .Y(_1656_) );
OAI22X1 OAI22X1_254 ( .A(_1654_), .B(_1547__bF_buf3), .C(_1601__bF_buf4), .D(_1656_), .Y(_2__21_) );
OAI22X1 OAI22X1_255 ( .A(_4499__bF_buf3), .B(_10559_), .C(_4500_), .D(_1510_), .Y(_1657_) );
NOR2X1 NOR2X1_1128 ( .A(_1657_), .B(_1630__bF_buf2), .Y(_1658_) );
OAI22X1 OAI22X1_256 ( .A(_9269_), .B(_1547__bF_buf2), .C(_1601__bF_buf3), .D(_1658_), .Y(_2__22_) );
INVX1 INVX1_1056 ( .A(decoded_imm_23_), .Y(_1659_) );
INVX1 INVX1_1057 ( .A(mem_rdata_q_23_), .Y(_1660_) );
OAI22X1 OAI22X1_257 ( .A(_4499__bF_buf2), .B(_10579_), .C(_4500_), .D(_1660_), .Y(_1661_) );
NOR2X1 NOR2X1_1129 ( .A(_1661_), .B(_1630__bF_buf1), .Y(_1662_) );
OAI22X1 OAI22X1_258 ( .A(_1659_), .B(_1547__bF_buf1), .C(_1601__bF_buf2), .D(_1662_), .Y(_2__23_) );
OAI21X1 OAI21X1_2522 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_24_), .Y(_1663_) );
OAI21X1 OAI21X1_2523 ( .A(_4499__bF_buf1), .B(_10612_), .C(_1663_), .Y(_1664_) );
NOR2X1 NOR2X1_1130 ( .A(_1664_), .B(_1630__bF_buf0), .Y(_1665_) );
OAI22X1 OAI22X1_259 ( .A(_9440_), .B(_1547__bF_buf0), .C(_1601__bF_buf1), .D(_1665_), .Y(_2__24_) );
OAI21X1 OAI21X1_2524 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_25_), .Y(_1666_) );
OAI21X1 OAI21X1_2525 ( .A(_4499__bF_buf0), .B(_10632_), .C(_1666_), .Y(_1667_) );
NOR2X1 NOR2X1_1131 ( .A(_1667_), .B(_1630__bF_buf3), .Y(_1668_) );
OAI22X1 OAI22X1_260 ( .A(_9520_), .B(_1547__bF_buf5), .C(_1601__bF_buf0), .D(_1668_), .Y(_2__25_) );
OAI21X1 OAI21X1_2526 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_26_), .Y(_1669_) );
OAI21X1 OAI21X1_2527 ( .A(_4499__bF_buf5), .B(_10652_), .C(_1669_), .Y(_1670_) );
NOR2X1 NOR2X1_1132 ( .A(_1670_), .B(_1630__bF_buf2), .Y(_1671_) );
OAI22X1 OAI22X1_261 ( .A(_9607_), .B(_1547__bF_buf4), .C(_1601__bF_buf4), .D(_1671_), .Y(_2__26_) );
INVX1 INVX1_1058 ( .A(mem_rdata_q_27_), .Y(_1672_) );
OAI22X1 OAI22X1_262 ( .A(_4499__bF_buf4), .B(_10670_), .C(_4500_), .D(_1672_), .Y(_1673_) );
NOR2X1 NOR2X1_1133 ( .A(_1673_), .B(_1630__bF_buf1), .Y(_1674_) );
OAI22X1 OAI22X1_263 ( .A(_9683_), .B(_1547__bF_buf3), .C(_1601__bF_buf3), .D(_1674_), .Y(_2__27_) );
OAI21X1 OAI21X1_2528 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_28_), .Y(_1675_) );
OAI21X1 OAI21X1_2529 ( .A(_4499__bF_buf3), .B(_10700_), .C(_1675_), .Y(_1676_) );
NOR2X1 NOR2X1_1134 ( .A(_1676_), .B(_1630__bF_buf0), .Y(_1677_) );
OAI22X1 OAI22X1_264 ( .A(_9770_), .B(_1547__bF_buf2), .C(_1601__bF_buf2), .D(_1677_), .Y(_2__28_) );
OAI21X1 OAI21X1_2530 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_29_), .Y(_1678_) );
OAI21X1 OAI21X1_2531 ( .A(_4499__bF_buf2), .B(_10716_), .C(_1678_), .Y(_1679_) );
NOR2X1 NOR2X1_1135 ( .A(_1679_), .B(_1630__bF_buf3), .Y(_1680_) );
OAI22X1 OAI22X1_265 ( .A(_9859_), .B(_1547__bF_buf1), .C(_1601__bF_buf1), .D(_1680_), .Y(_2__29_) );
INVX1 INVX1_1059 ( .A(mem_rdata_q_30_), .Y(_1681_) );
OAI22X1 OAI22X1_266 ( .A(_4499__bF_buf1), .B(_1528_), .C(_4500_), .D(_1681_), .Y(_1682_) );
NOR2X1 NOR2X1_1136 ( .A(_1682_), .B(_1630__bF_buf2), .Y(_1683_) );
OAI22X1 OAI22X1_267 ( .A(_9943_), .B(_1547__bF_buf0), .C(_1601__bF_buf0), .D(_1683_), .Y(_2__30_) );
OAI21X1 OAI21X1_2532 ( .A(_4605__bF_buf3), .B(decoder_pseudo_trigger_bF_buf1), .C(decoded_imm_31_), .Y(_1684_) );
OAI21X1 OAI21X1_2533 ( .A(instr_lui), .B(instr_auipc), .C(mem_rdata_q_31_), .Y(_1685_) );
OAI21X1 OAI21X1_2534 ( .A(_4499__bF_buf0), .B(_1169_), .C(_1685_), .Y(_1686_) );
NOR2X1 NOR2X1_1137 ( .A(_1686_), .B(_1630__bF_buf1), .Y(_1687_) );
OAI21X1 OAI21X1_2535 ( .A(_1601__bF_buf4), .B(_1687_), .C(_1684_), .Y(_2__31_) );
OAI21X1 OAI21X1_2536 ( .A(_5362__bF_buf0), .B(_4985__bF_buf8), .C(_1534_), .Y(_6__0_) );
OAI21X1 OAI21X1_2537 ( .A(_5349__bF_buf6), .B(_4985__bF_buf7), .C(_1509_), .Y(_6__1_) );
OAI21X1 OAI21X1_2538 ( .A(_5358__bF_buf11), .B(_4985__bF_buf6), .C(_1512_), .Y(_6__2_) );
OAI21X1 OAI21X1_2539 ( .A(_5348__bF_buf1), .B(_4985__bF_buf5), .C(_1515_), .Y(_6__3_) );
OAI21X1 OAI21X1_2540 ( .A(_5347_), .B(_4985__bF_buf4), .C(_1531_), .Y(_6__4_) );
NAND2X1 NAND2X1_849 ( .A(mem_rdata_latched_12_), .B(_4985__bF_buf3), .Y(_1688_) );
OAI21X1 OAI21X1_2541 ( .A(_10347_), .B(_4985__bF_buf2), .C(_1688_), .Y(_3__12_) );
NAND2X1 NAND2X1_850 ( .A(mem_rdata_latched_13_), .B(_4985__bF_buf1), .Y(_1689_) );
OAI21X1 OAI21X1_2542 ( .A(_10360_), .B(_4985__bF_buf0), .C(_1689_), .Y(_3__13_) );
NAND2X1 NAND2X1_851 ( .A(mem_rdata_latched_14_), .B(_4985__bF_buf8), .Y(_1690_) );
OAI21X1 OAI21X1_2543 ( .A(_10382_), .B(_4985__bF_buf7), .C(_1690_), .Y(_3__14_) );
OAI21X1 OAI21X1_2544 ( .A(_10397_), .B(_4985__bF_buf6), .C(_1537_), .Y(_3__15_) );
OAI21X1 OAI21X1_2545 ( .A(_10433_), .B(_4985__bF_buf5), .C(_1540_), .Y(_3__16_) );
OAI21X1 OAI21X1_2546 ( .A(_10454_), .B(_4985__bF_buf4), .C(_1543_), .Y(_3__17_) );
OAI21X1 OAI21X1_2547 ( .A(_10470_), .B(_4985__bF_buf3), .C(_1546_), .Y(_3__18_) );
OAI21X1 OAI21X1_2548 ( .A(_10490_), .B(_4985__bF_buf2), .C(_1497_), .Y(_3__19_) );
NAND2X1 NAND2X1_852 ( .A(mem_rdata[7]), .B(_4542_), .Y(_1691_) );
OAI21X1 OAI21X1_2549 ( .A(_1594_), .B(_4542_), .C(_1691_), .Y(mem_rdata_latched_7_) );
NAND2X1 NAND2X1_853 ( .A(mem_rdata_latched_7_), .B(_4985__bF_buf1), .Y(_1692_) );
OAI21X1 OAI21X1_2550 ( .A(_5736_), .B(_4985__bF_buf0), .C(_1692_), .Y(_4__0_) );
INVX1 INVX1_1060 ( .A(mem_rdata[8]), .Y(_1693_) );
NAND2X1 NAND2X1_854 ( .A(mem_rdata_q_8_), .B(_4439__bF_buf3), .Y(_1694_) );
OAI21X1 OAI21X1_2551 ( .A(_1693_), .B(_4439__bF_buf2), .C(_1694_), .Y(mem_rdata_latched_8_) );
NAND2X1 NAND2X1_855 ( .A(mem_rdata_latched_8_), .B(_4985__bF_buf8), .Y(_1695_) );
OAI21X1 OAI21X1_2552 ( .A(_5740_), .B(_4985__bF_buf7), .C(_1695_), .Y(_4__1_) );
INVX1 INVX1_1061 ( .A(mem_rdata[9]), .Y(_1696_) );
NAND2X1 NAND2X1_856 ( .A(mem_rdata_q_9_), .B(_4439__bF_buf1), .Y(_1697_) );
OAI21X1 OAI21X1_2553 ( .A(_1696_), .B(_4439__bF_buf0), .C(_1697_), .Y(mem_rdata_latched_9_) );
NAND2X1 NAND2X1_857 ( .A(mem_rdata_latched_9_), .B(_4985__bF_buf6), .Y(_1698_) );
OAI21X1 OAI21X1_2554 ( .A(_5741_), .B(_4985__bF_buf5), .C(_1698_), .Y(_4__2_) );
INVX1 INVX1_1062 ( .A(mem_rdata[10]), .Y(_1699_) );
NAND2X1 NAND2X1_858 ( .A(mem_rdata_q_10_), .B(_4439__bF_buf6), .Y(_1700_) );
OAI21X1 OAI21X1_2555 ( .A(_1699_), .B(_4439__bF_buf5), .C(_1700_), .Y(mem_rdata_latched_10_) );
NAND2X1 NAND2X1_859 ( .A(mem_rdata_latched_10_), .B(_4985__bF_buf4), .Y(_1701_) );
OAI21X1 OAI21X1_2556 ( .A(_5742_), .B(_4985__bF_buf3), .C(_1701_), .Y(_4__3_) );
INVX1 INVX1_1063 ( .A(mem_rdata[11]), .Y(_1702_) );
NAND2X1 NAND2X1_860 ( .A(mem_rdata_q_11_), .B(_4439__bF_buf4), .Y(_1703_) );
OAI21X1 OAI21X1_2557 ( .A(_1702_), .B(_4439__bF_buf3), .C(_1703_), .Y(mem_rdata_latched_11_) );
NAND2X1 NAND2X1_861 ( .A(mem_rdata_latched_11_), .B(_4985__bF_buf2), .Y(_1704_) );
OAI21X1 OAI21X1_2558 ( .A(_5744_), .B(_4985__bF_buf1), .C(_1704_), .Y(_4__4_) );
OAI21X1 OAI21X1_2559 ( .A(_4605__bF_buf2), .B(decoder_pseudo_trigger_bF_buf0), .C(instr_rdinstrh), .Y(_1705_) );
NOR2X1 NOR2X1_1138 ( .A(mem_rdata_q_2_), .B(mem_rdata_q_19_), .Y(_1706_) );
NAND3X1 NAND3X1_87 ( .A(_1636_), .B(_1538_), .C(_1706_), .Y(_1707_) );
AND2X2 AND2X2_199 ( .A(mem_rdata_q_5_), .B(mem_rdata_q_6_), .Y(_1708_) );
NAND3X1 NAND3X1_88 ( .A(_4541_), .B(mem_rdata_q_4_), .C(_1708_), .Y(_1709_) );
NOR2X1 NOR2X1_1139 ( .A(_1707_), .B(_1709_), .Y(_1710_) );
NOR2X1 NOR2X1_1140 ( .A(mem_rdata_q_12_), .B(_1631_), .Y(_1711_) );
INVX1 INVX1_1064 ( .A(_1711_), .Y(_1712_) );
NOR2X1 NOR2X1_1141 ( .A(mem_rdata_q_14_), .B(_1712_), .Y(_1713_) );
INVX1 INVX1_1065 ( .A(_1713_), .Y(_1714_) );
NOR2X1 NOR2X1_1142 ( .A(mem_rdata_q_17_), .B(mem_rdata_q_18_), .Y(_1715_) );
NAND3X1 NAND3X1_89 ( .A(mem_rdata_q_0_), .B(mem_rdata_q_1_), .C(_1715_), .Y(_1716_) );
NOR2X1 NOR2X1_1143 ( .A(_1716_), .B(_1714_), .Y(_1717_) );
NAND2X1 NAND2X1_862 ( .A(_1710_), .B(_1717_), .Y(_1718_) );
NAND2X1 NAND2X1_863 ( .A(mem_rdata_q_30_), .B(mem_rdata_q_31_), .Y(_1719_) );
NOR3X1 NOR3X1_7 ( .A(mem_rdata_q_28_), .B(mem_rdata_q_29_), .C(_1719_), .Y(_1720_) );
INVX1 INVX1_1066 ( .A(_1720_), .Y(_1721_) );
NOR2X1 NOR2X1_1144 ( .A(mem_rdata_q_25_), .B(mem_rdata_q_24_), .Y(_1722_) );
NOR2X1 NOR2X1_1145 ( .A(mem_rdata_q_26_), .B(_1672_), .Y(_1723_) );
NAND2X1 NAND2X1_864 ( .A(_1722_), .B(_1723_), .Y(_1724_) );
NOR2X1 NOR2X1_1146 ( .A(_1724_), .B(_1721_), .Y(_1725_) );
NAND2X1 NAND2X1_865 ( .A(_1510_), .B(_1660_), .Y(_1726_) );
NOR2X1 NOR2X1_1147 ( .A(mem_rdata_q_20_), .B(_1507_), .Y(_1727_) );
NAND2X1 NAND2X1_866 ( .A(_1547__bF_buf5), .B(_1727_), .Y(_1728_) );
NOR2X1 NOR2X1_1148 ( .A(_1726_), .B(_1728_), .Y(_1729_) );
NAND2X1 NAND2X1_867 ( .A(_1729_), .B(_1725_), .Y(_1730_) );
OAI21X1 OAI21X1_2560 ( .A(_1718_), .B(_1730_), .C(_1705_), .Y(_33_) );
INVX1 INVX1_1067 ( .A(_1718_), .Y(_1731_) );
NAND2X1 NAND2X1_868 ( .A(_1569_), .B(_1722_), .Y(_1732_) );
NOR2X1 NOR2X1_1149 ( .A(_1732_), .B(_1721_), .Y(_1733_) );
NAND3X1 NAND3X1_90 ( .A(_1729_), .B(_1733_), .C(_1731_), .Y(_1734_) );
OAI21X1 OAI21X1_2561 ( .A(_4529_), .B(_1547__bF_buf4), .C(_1734_), .Y(_32_) );
INVX1 INVX1_1068 ( .A(instr_rdcycleh_bF_buf2), .Y(_1735_) );
INVX1 INVX1_1069 ( .A(_1725_), .Y(_1736_) );
NAND2X1 NAND2X1_869 ( .A(_1507_), .B(_1547__bF_buf3), .Y(_1737_) );
NOR2X1 NOR2X1_1150 ( .A(_1726_), .B(_1737_), .Y(_1738_) );
NAND2X1 NAND2X1_870 ( .A(_1738_), .B(_1731_), .Y(_1739_) );
OAI22X1 OAI22X1_268 ( .A(_1735_), .B(_1547__bF_buf2), .C(_1739_), .D(_1736_), .Y(_31_) );
INVX1 INVX1_1070 ( .A(_1733_), .Y(_1740_) );
OAI21X1 OAI21X1_2562 ( .A(_4605__bF_buf1), .B(decoder_pseudo_trigger_bF_buf3), .C(instr_rdcycle_bF_buf3), .Y(_1741_) );
OAI21X1 OAI21X1_2563 ( .A(_1739_), .B(_1740_), .C(_1741_), .Y(_30_) );
NOR2X1 NOR2X1_1151 ( .A(_1575_), .B(_1578_), .Y(_1742_) );
NAND2X1 NAND2X1_871 ( .A(is_alu_reg_imm), .B(_1742_), .Y(_1743_) );
NOR2X1 NOR2X1_1152 ( .A(_1681_), .B(_1566__bF_buf0), .Y(_1744_) );
NAND2X1 NAND2X1_872 ( .A(_1574_), .B(_1744_), .Y(_1745_) );
OAI22X1 OAI22X1_269 ( .A(_4517_), .B(_1547__bF_buf1), .C(_1743_), .D(_1745_), .Y(_43_) );
NAND2X1 NAND2X1_873 ( .A(_1681_), .B(_1574_), .Y(_1746_) );
NOR2X1 NOR2X1_1153 ( .A(_1566__bF_buf3), .B(_1746_), .Y(_1747_) );
INVX1 INVX1_1071 ( .A(_1747_), .Y(_1748_) );
OAI22X1 OAI22X1_270 ( .A(_4516_), .B(_1547__bF_buf0), .C(_1748_), .D(_1743_), .Y(_45_) );
OAI21X1 OAI21X1_2564 ( .A(_4605__bF_buf0), .B(decoder_pseudo_trigger_bF_buf2), .C(instr_slli), .Y(_1749_) );
NOR2X1 NOR2X1_1154 ( .A(mem_rdata_q_14_), .B(_1578_), .Y(_1750_) );
NAND2X1 NAND2X1_874 ( .A(_1584_), .B(_1750_), .Y(_1751_) );
OAI21X1 OAI21X1_2565 ( .A(_1751_), .B(_1746_), .C(_1749_), .Y(_37_) );
NAND2X1 NAND2X1_875 ( .A(is_sb_sh_sw), .B(_1547__bF_buf5), .Y(_1752_) );
OAI21X1 OAI21X1_2566 ( .A(_4605__bF_buf5), .B(decoder_pseudo_trigger_bF_buf1), .C(instr_sw), .Y(_1753_) );
OAI21X1 OAI21X1_2567 ( .A(_1714_), .B(_1752_), .C(_1753_), .Y(_47_) );
INVX1 INVX1_1072 ( .A(_1750_), .Y(_1754_) );
OAI21X1 OAI21X1_2568 ( .A(_4605__bF_buf4), .B(decoder_pseudo_trigger_bF_buf0), .C(instr_sh), .Y(_1755_) );
OAI21X1 OAI21X1_2569 ( .A(_1754_), .B(_1752_), .C(_1755_), .Y(_35_) );
NAND2X1 NAND2X1_876 ( .A(_1576_), .B(_1631_), .Y(_1756_) );
NOR2X1 NOR2X1_1155 ( .A(mem_rdata_q_14_), .B(_1756_), .Y(_1757_) );
INVX1 INVX1_1073 ( .A(_1757_), .Y(_1758_) );
OAI21X1 OAI21X1_2570 ( .A(_4605__bF_buf3), .B(decoder_pseudo_trigger_bF_buf3), .C(instr_sb), .Y(_1759_) );
OAI21X1 OAI21X1_2571 ( .A(_1758_), .B(_1752_), .C(_1759_), .Y(_34_) );
INVX1 INVX1_1074 ( .A(_1742_), .Y(_1760_) );
NAND2X1 NAND2X1_877 ( .A(is_lb_lh_lw_lbu_lhu), .B(_1547__bF_buf4), .Y(_1761_) );
OAI21X1 OAI21X1_2572 ( .A(_4605__bF_buf2), .B(decoder_pseudo_trigger_bF_buf2), .C(instr_lhu), .Y(_1762_) );
OAI21X1 OAI21X1_2573 ( .A(_1760_), .B(_1761_), .C(_1762_), .Y(_25_) );
OR2X2 OR2X2_39 ( .A(_1756_), .B(_1575_), .Y(_1763_) );
OAI21X1 OAI21X1_2574 ( .A(_4605__bF_buf1), .B(decoder_pseudo_trigger_bF_buf1), .C(instr_lbu), .Y(_1764_) );
OAI21X1 OAI21X1_2575 ( .A(_1763_), .B(_1761_), .C(_1764_), .Y(_23_) );
OAI22X1 OAI22X1_271 ( .A(_4521_), .B(_1547__bF_buf3), .C(_1714_), .D(_1761_), .Y(_27_) );
OAI21X1 OAI21X1_2576 ( .A(_4605__bF_buf0), .B(decoder_pseudo_trigger_bF_buf0), .C(instr_lh), .Y(_1765_) );
OAI21X1 OAI21X1_2577 ( .A(_1754_), .B(_1761_), .C(_1765_), .Y(_24_) );
OAI21X1 OAI21X1_2578 ( .A(_4605__bF_buf5), .B(decoder_pseudo_trigger_bF_buf3), .C(instr_lb), .Y(_1766_) );
OAI21X1 OAI21X1_2579 ( .A(_1758_), .B(_1761_), .C(_1766_), .Y(_22_) );
NAND2X1 NAND2X1_878 ( .A(mem_rdata_latched_2_), .B(_1558_), .Y(_1767_) );
NOR2X1 NOR2X1_1156 ( .A(mem_rdata_latched_3_), .B(_1767_), .Y(_1768_) );
AND2X2 AND2X2_200 ( .A(_1581_), .B(mem_rdata_latched_6_), .Y(_1769_) );
OR2X2 OR2X2_40 ( .A(mem_rdata_latched_12_), .B(mem_rdata_latched_13_), .Y(_1770_) );
NOR2X1 NOR2X1_1157 ( .A(mem_rdata_latched_14_), .B(_1770_), .Y(_1771_) );
NAND3X1 NAND3X1_91 ( .A(_1768_), .B(_1771_), .C(_1769_), .Y(_1772_) );
OAI21X1 OAI21X1_2580 ( .A(_4588_), .B(_4984_), .C(instr_jalr), .Y(_1773_) );
OAI21X1 OAI21X1_2581 ( .A(_1772_), .B(_1587_), .C(_1773_), .Y(_21_) );
INVX1 INVX1_1075 ( .A(_1767_), .Y(_1774_) );
NAND3X1 NAND3X1_92 ( .A(mem_rdata_latched_3_), .B(_1774_), .C(_1769_), .Y(_1775_) );
OAI21X1 OAI21X1_2582 ( .A(_4588_), .B(_4984_), .C(instr_jal_bF_buf1), .Y(_1776_) );
OAI21X1 OAI21X1_2583 ( .A(_1775_), .B(_1587_), .C(_1776_), .Y(_20_) );
NAND2X1 NAND2X1_879 ( .A(_1564_), .B(_1768_), .Y(_1777_) );
OAI21X1 OAI21X1_2584 ( .A(_4588_), .B(_4984_), .C(instr_auipc), .Y(_1778_) );
OAI21X1 OAI21X1_2585 ( .A(_1777_), .B(_1587_), .C(_1778_), .Y(_13_) );
NAND2X1 NAND2X1_880 ( .A(_1556_), .B(_1768_), .Y(_1779_) );
OAI21X1 OAI21X1_2586 ( .A(_4588_), .B(_4984_), .C(instr_lui), .Y(_1780_) );
OAI21X1 OAI21X1_2587 ( .A(_1779_), .B(_1587_), .C(_1780_), .Y(_26_) );
NAND2X1 NAND2X1_881 ( .A(resetn_bF_buf2), .B(_10736_), .Y(_1781_) );
NOR2X1 NOR2X1_1158 ( .A(_10736_), .B(_4426__bF_buf3), .Y(_1782_) );
NOR2X1 NOR2X1_1159 ( .A(mem_do_rdata), .B(_4621__bF_buf3), .Y(_1783_) );
NAND2X1 NAND2X1_882 ( .A(_4435_), .B(_4438_), .Y(_1784_) );
NOR2X1 NOR2X1_1160 ( .A(_1784_), .B(_1783_), .Y(_1785_) );
NAND2X1 NAND2X1_883 ( .A(mem_state_0_), .B(_4432_), .Y(_1786_) );
NOR2X1 NOR2X1_1161 ( .A(_4439__bF_buf2), .B(_4436_), .Y(_1787_) );
NAND2X1 NAND2X1_884 ( .A(_4984_), .B(_4434_), .Y(_1788_) );
OAI21X1 OAI21X1_2588 ( .A(_1786_), .B(_1787_), .C(_1788_), .Y(_1789_) );
OAI21X1 OAI21X1_2589 ( .A(_1785_), .B(_1789_), .C(_1782_), .Y(_1790_) );
OAI21X1 OAI21X1_2590 ( .A(_4433_), .B(_1781_), .C(_1790_), .Y(_76__0_) );
NOR2X1 NOR2X1_1162 ( .A(_4435_), .B(_4619_), .Y(_1791_) );
NAND2X1 NAND2X1_885 ( .A(_4436_), .B(_4542_), .Y(_1792_) );
NOR2X1 NOR2X1_1163 ( .A(mem_state_0_), .B(_4432_), .Y(_1793_) );
AOI22X1 AOI22X1_112 ( .A(_1793_), .B(_4439__bF_buf1), .C(_4984_), .D(_4434_), .Y(_1794_) );
OAI21X1 OAI21X1_2591 ( .A(_1786_), .B(_1792_), .C(_1794_), .Y(_1795_) );
OAI21X1 OAI21X1_2592 ( .A(_1795_), .B(_1791_), .C(_1782_), .Y(_1796_) );
OAI21X1 OAI21X1_2593 ( .A(_4432_), .B(_1781_), .C(_1796_), .Y(_76__1_) );
INVX1 INVX1_1076 ( .A(mem_wordsize_2_), .Y(_1797_) );
OAI21X1 OAI21X1_2594 ( .A(_1797_), .B(_10734__1_), .C(_4425_), .Y(_1798_) );
INVX1 INVX1_1077 ( .A(_1798_), .Y(_1799_) );
OAI21X1 OAI21X1_2595 ( .A(_10734__1_), .B(_10734__0_), .C(_1799_), .Y(_10730__0_) );
OAI21X1 OAI21X1_2596 ( .A(_4426__bF_buf2), .B(_10736_), .C(_10733__0_), .Y(_1800_) );
OAI21X1 OAI21X1_2597 ( .A(_1783_), .B(_4619_), .C(_1782_), .Y(_1801_) );
NOR2X1 NOR2X1_1164 ( .A(_10729_), .B(_10727_), .Y(_1802_) );
AOI22X1 AOI22X1_113 ( .A(_10729_), .B(_10730__0_), .C(_1802_), .D(_10733__0_), .Y(_1803_) );
OAI21X1 OAI21X1_2598 ( .A(_1803_), .B(_1801_), .C(_1800_), .Y(_79__0_) );
OAI21X1 OAI21X1_2599 ( .A(_10734__1_), .B(_4491_), .C(_1799_), .Y(_10730__1_) );
OAI21X1 OAI21X1_2600 ( .A(_4426__bF_buf1), .B(_10736_), .C(_10733__1_), .Y(_1804_) );
AOI22X1 AOI22X1_114 ( .A(_10729_), .B(_10730__1_), .C(_1802_), .D(_10733__1_), .Y(_1805_) );
OAI21X1 OAI21X1_2601 ( .A(_1805_), .B(_1801_), .C(_1804_), .Y(_79__1_) );
NAND2X1 NAND2X1_886 ( .A(_10734__1_), .B(_4425_), .Y(_1806_) );
NOR2X1 NOR2X1_1165 ( .A(_1797_), .B(_4490_), .Y(_1807_) );
INVX1 INVX1_1078 ( .A(_1807_), .Y(_1808_) );
OAI21X1 OAI21X1_2602 ( .A(_1806_), .B(_10734__0_), .C(_1808_), .Y(_1809_) );
INVX1 INVX1_1079 ( .A(_1809_), .Y(_1810_) );
NAND2X1 NAND2X1_887 ( .A(_4425_), .B(_1810_), .Y(_10730__2_) );
OAI21X1 OAI21X1_2603 ( .A(_4426__bF_buf0), .B(_10736_), .C(_10733__2_), .Y(_1811_) );
AOI22X1 AOI22X1_115 ( .A(_1802_), .B(_10733__2_), .C(_10729_), .D(_10730__2_), .Y(_1812_) );
OAI21X1 OAI21X1_2604 ( .A(_1812_), .B(_1801_), .C(_1811_), .Y(_79__2_) );
OAI21X1 OAI21X1_2605 ( .A(mem_wordsize_2_), .B(_10734__0_), .C(_10734__1_), .Y(_1813_) );
NAND2X1 NAND2X1_888 ( .A(_4425_), .B(_1813_), .Y(_10730__3_) );
OAI21X1 OAI21X1_2606 ( .A(_4426__bF_buf11), .B(_10736_), .C(_10733__3_), .Y(_1814_) );
AOI22X1 AOI22X1_116 ( .A(_10729_), .B(_10730__3_), .C(_1802_), .D(_10733__3_), .Y(_1815_) );
OAI21X1 OAI21X1_2607 ( .A(_1815_), .B(_1801_), .C(_1814_), .Y(_79__3_) );
NOR2X1 NOR2X1_1166 ( .A(mem_wordsize_0_bF_buf1_), .B(mem_wordsize_2_), .Y(_1816_) );
INVX1 INVX1_1080 ( .A(_1816_), .Y(_1817_) );
NOR2X1 NOR2X1_1167 ( .A(_5142_), .B(_1817__bF_buf3), .Y(_1818_) );
AOI21X1 AOI21X1_861 ( .A(_10735__8_), .B(_1817__bF_buf2), .C(_1818_), .Y(_1819_) );
INVX1 INVX1_1081 ( .A(_1819_), .Y(_10728__8_) );
NOR2X1 NOR2X1_1168 ( .A(_5140__bF_buf2), .B(_1817__bF_buf1), .Y(_1820_) );
AOI21X1 AOI21X1_862 ( .A(_10735__9_), .B(_1817__bF_buf0), .C(_1820_), .Y(_1821_) );
INVX1 INVX1_1082 ( .A(_1821_), .Y(_10728__9_) );
NOR2X1 NOR2X1_1169 ( .A(_5131__bF_buf2), .B(_1817__bF_buf3), .Y(_1822_) );
AOI21X1 AOI21X1_863 ( .A(_10735__10_), .B(_1817__bF_buf2), .C(_1822_), .Y(_1823_) );
INVX1 INVX1_1083 ( .A(_1823_), .Y(_10728__10_) );
NOR2X1 NOR2X1_1170 ( .A(_5856__bF_buf3), .B(_1817__bF_buf1), .Y(_1824_) );
AOI21X1 AOI21X1_864 ( .A(_10735__11_), .B(_1817__bF_buf0), .C(_1824_), .Y(_1825_) );
INVX1 INVX1_1084 ( .A(_1825_), .Y(_10728__11_) );
NOR2X1 NOR2X1_1171 ( .A(_5859__bF_buf3), .B(_1817__bF_buf3), .Y(_1826_) );
AOI21X1 AOI21X1_865 ( .A(_10735__12_), .B(_1817__bF_buf2), .C(_1826_), .Y(_1827_) );
INVX1 INVX1_1085 ( .A(_1827_), .Y(_10728__12_) );
NOR2X1 NOR2X1_1172 ( .A(_5862_), .B(_1817__bF_buf1), .Y(_1828_) );
AOI21X1 AOI21X1_866 ( .A(_10735__13_), .B(_1817__bF_buf0), .C(_1828_), .Y(_1829_) );
INVX1 INVX1_1086 ( .A(_1829_), .Y(_10728__13_) );
NOR2X1 NOR2X1_1173 ( .A(_5926_), .B(_1817__bF_buf3), .Y(_1830_) );
AOI21X1 AOI21X1_867 ( .A(_10735__14_), .B(_1817__bF_buf2), .C(_1830_), .Y(_1831_) );
INVX1 INVX1_1087 ( .A(_1831_), .Y(_10728__14_) );
NOR2X1 NOR2X1_1174 ( .A(_5990_), .B(_1817__bF_buf1), .Y(_1832_) );
AOI21X1 AOI21X1_868 ( .A(_10735__15_), .B(_1817__bF_buf0), .C(_1832_), .Y(_1833_) );
INVX1 INVX1_1088 ( .A(_1833_), .Y(_10728__15_) );
NOR2X1 NOR2X1_1175 ( .A(mem_wordsize_2_), .B(_4425_), .Y(_1834_) );
INVX1 INVX1_1089 ( .A(_1834_), .Y(_1835_) );
AOI22X1 AOI22X1_117 ( .A(mem_wordsize_0_bF_buf0_), .B(_10735__16_), .C(_1835_), .D(_10728__0_bF_buf4_), .Y(_1836_) );
INVX1 INVX1_1090 ( .A(_1836_), .Y(_10728__16_) );
AOI22X1 AOI22X1_118 ( .A(mem_wordsize_0_bF_buf3_), .B(_10735__17_), .C(_1835_), .D(_10728__1_bF_buf1_), .Y(_1837_) );
INVX1 INVX1_1091 ( .A(_1837_), .Y(_10728__17_) );
AOI22X1 AOI22X1_119 ( .A(mem_wordsize_0_bF_buf2_), .B(_10735__18_), .C(_1835_), .D(_10728__2_bF_buf2_), .Y(_1838_) );
INVX1 INVX1_1092 ( .A(_1838_), .Y(_10728__18_) );
AOI22X1 AOI22X1_120 ( .A(mem_wordsize_0_bF_buf1_), .B(_10735__19_), .C(_1835_), .D(_10728__3_bF_buf0_), .Y(_1839_) );
INVX1 INVX1_1093 ( .A(_1839_), .Y(_10728__19_) );
AOI22X1 AOI22X1_121 ( .A(mem_wordsize_0_bF_buf0_), .B(_10735__20_), .C(_1835_), .D(_10728__4_bF_buf0_), .Y(_1840_) );
INVX1 INVX1_1094 ( .A(_1840_), .Y(_10728__20_) );
AOI22X1 AOI22X1_122 ( .A(mem_wordsize_0_bF_buf3_), .B(_10735__21_), .C(_1835_), .D(_10728__5_), .Y(_1841_) );
INVX1 INVX1_1095 ( .A(_1841_), .Y(_10728__21_) );
AOI22X1 AOI22X1_123 ( .A(mem_wordsize_0_bF_buf2_), .B(_10735__22_), .C(_1835_), .D(_10728__6_), .Y(_1842_) );
INVX1 INVX1_1096 ( .A(_1842_), .Y(_10728__22_) );
AOI22X1 AOI22X1_124 ( .A(mem_wordsize_0_bF_buf1_), .B(_10735__23_), .C(_1835_), .D(_10728__7_), .Y(_1843_) );
INVX1 INVX1_1097 ( .A(_1843_), .Y(_10728__23_) );
AOI21X1 AOI21X1_869 ( .A(mem_wordsize_0_bF_buf0_), .B(_10735__24_), .C(_1818_), .Y(_1844_) );
OAI21X1 OAI21X1_2608 ( .A(_1797_), .B(_6051_), .C(_1844_), .Y(_10728__24_) );
AOI21X1 AOI21X1_870 ( .A(mem_wordsize_0_bF_buf3_), .B(_10735__25_), .C(_1820_), .Y(_1845_) );
OAI21X1 OAI21X1_2609 ( .A(_1797_), .B(_5108_), .C(_1845_), .Y(_10728__25_) );
AOI21X1 AOI21X1_871 ( .A(mem_wordsize_0_bF_buf2_), .B(_10735__26_), .C(_1822_), .Y(_1846_) );
OAI21X1 OAI21X1_2610 ( .A(_1797_), .B(_5122_), .C(_1846_), .Y(_10728__26_) );
AOI21X1 AOI21X1_872 ( .A(mem_wordsize_0_bF_buf1_), .B(_10735__27_), .C(_1824_), .Y(_1847_) );
OAI21X1 OAI21X1_2611 ( .A(_1797_), .B(_5118_), .C(_1847_), .Y(_10728__27_) );
AOI22X1 AOI22X1_125 ( .A(mem_wordsize_0_bF_buf0_), .B(_10735__28_), .C(mem_wordsize_2_), .D(_10735__12_), .Y(_1848_) );
OAI21X1 OAI21X1_2612 ( .A(_1817__bF_buf3), .B(_5859__bF_buf2), .C(_1848_), .Y(_10728__28_) );
AOI22X1 AOI22X1_126 ( .A(mem_wordsize_0_bF_buf3_), .B(_10735__29_), .C(mem_wordsize_2_), .D(_10735__13_), .Y(_1849_) );
OAI21X1 OAI21X1_2613 ( .A(_1817__bF_buf2), .B(_5862_), .C(_1849_), .Y(_10728__29_) );
AOI22X1 AOI22X1_127 ( .A(mem_wordsize_0_bF_buf2_), .B(_10735__30_), .C(mem_wordsize_2_), .D(_10735__14_), .Y(_1850_) );
OAI21X1 OAI21X1_2614 ( .A(_1817__bF_buf1), .B(_5926_), .C(_1850_), .Y(_10728__30_) );
AOI21X1 AOI21X1_873 ( .A(mem_wordsize_0_bF_buf1_), .B(_10735__31_), .C(_1832_), .Y(_1851_) );
OAI21X1 OAI21X1_2615 ( .A(_1797_), .B(_5088_), .C(_1851_), .Y(_10728__31_) );
INVX1 INVX1_1098 ( .A(_10732__0_), .Y(_1852_) );
NAND2X1 NAND2X1_889 ( .A(_1782_), .B(_1791_), .Y(_1853_) );
MUX2X1 MUX2X1_233 ( .A(_1852_), .B(_5142_), .S(_1853__bF_buf5), .Y(_78__0_) );
INVX1 INVX1_1099 ( .A(_10732__1_), .Y(_1854_) );
MUX2X1 MUX2X1_234 ( .A(_1854_), .B(_5140__bF_buf1), .S(_1853__bF_buf4), .Y(_78__1_) );
INVX1 INVX1_1100 ( .A(_10732__2_), .Y(_1855_) );
MUX2X1 MUX2X1_235 ( .A(_1855_), .B(_5131__bF_buf1), .S(_1853__bF_buf3), .Y(_78__2_) );
INVX1 INVX1_1101 ( .A(_10732__3_), .Y(_1856_) );
MUX2X1 MUX2X1_236 ( .A(_1856_), .B(_5856__bF_buf2), .S(_1853__bF_buf2), .Y(_78__3_) );
INVX1 INVX1_1102 ( .A(_10732__4_), .Y(_1857_) );
MUX2X1 MUX2X1_237 ( .A(_1857_), .B(_5859__bF_buf1), .S(_1853__bF_buf1), .Y(_78__4_) );
INVX1 INVX1_1103 ( .A(_10732__5_), .Y(_1858_) );
MUX2X1 MUX2X1_238 ( .A(_1858_), .B(_5862_), .S(_1853__bF_buf0), .Y(_78__5_) );
INVX1 INVX1_1104 ( .A(_10732__6_), .Y(_1859_) );
MUX2X1 MUX2X1_239 ( .A(_1859_), .B(_5926_), .S(_1853__bF_buf5), .Y(_78__6_) );
INVX1 INVX1_1105 ( .A(_10732__7_), .Y(_1860_) );
MUX2X1 MUX2X1_240 ( .A(_1860_), .B(_5990_), .S(_1853__bF_buf4), .Y(_78__7_) );
INVX1 INVX1_1106 ( .A(_10732__8_), .Y(_1861_) );
MUX2X1 MUX2X1_241 ( .A(_1861_), .B(_1819_), .S(_1853__bF_buf3), .Y(_78__8_) );
INVX1 INVX1_1107 ( .A(_10732__9_), .Y(_1862_) );
MUX2X1 MUX2X1_242 ( .A(_1862_), .B(_1821_), .S(_1853__bF_buf2), .Y(_78__9_) );
INVX1 INVX1_1108 ( .A(_10732__10_), .Y(_1863_) );
MUX2X1 MUX2X1_243 ( .A(_1863_), .B(_1823_), .S(_1853__bF_buf1), .Y(_78__10_) );
INVX1 INVX1_1109 ( .A(_10732__11_), .Y(_1864_) );
MUX2X1 MUX2X1_244 ( .A(_1864_), .B(_1825_), .S(_1853__bF_buf0), .Y(_78__11_) );
INVX1 INVX1_1110 ( .A(_10732__12_), .Y(_1865_) );
MUX2X1 MUX2X1_245 ( .A(_1865_), .B(_1827_), .S(_1853__bF_buf5), .Y(_78__12_) );
INVX1 INVX1_1111 ( .A(_10732__13_), .Y(_1866_) );
MUX2X1 MUX2X1_246 ( .A(_1866_), .B(_1829_), .S(_1853__bF_buf4), .Y(_78__13_) );
INVX1 INVX1_1112 ( .A(_10732__14_), .Y(_1867_) );
MUX2X1 MUX2X1_247 ( .A(_1867_), .B(_1831_), .S(_1853__bF_buf3), .Y(_78__14_) );
INVX1 INVX1_1113 ( .A(_10732__15_), .Y(_1868_) );
MUX2X1 MUX2X1_248 ( .A(_1868_), .B(_1833_), .S(_1853__bF_buf2), .Y(_78__15_) );
INVX1 INVX1_1114 ( .A(_10732__16_), .Y(_1869_) );
MUX2X1 MUX2X1_249 ( .A(_1869_), .B(_1836_), .S(_1853__bF_buf1), .Y(_78__16_) );
INVX1 INVX1_1115 ( .A(_10732__17_), .Y(_1870_) );
MUX2X1 MUX2X1_250 ( .A(_1870_), .B(_1837_), .S(_1853__bF_buf0), .Y(_78__17_) );
INVX1 INVX1_1116 ( .A(_10732__18_), .Y(_1871_) );
MUX2X1 MUX2X1_251 ( .A(_1871_), .B(_1838_), .S(_1853__bF_buf5), .Y(_78__18_) );
INVX1 INVX1_1117 ( .A(_10732__19_), .Y(_1872_) );
MUX2X1 MUX2X1_252 ( .A(_1872_), .B(_1839_), .S(_1853__bF_buf4), .Y(_78__19_) );
INVX1 INVX1_1118 ( .A(_10732__20_), .Y(_1873_) );
MUX2X1 MUX2X1_253 ( .A(_1873_), .B(_1840_), .S(_1853__bF_buf3), .Y(_78__20_) );
INVX1 INVX1_1119 ( .A(_10732__21_), .Y(_1874_) );
MUX2X1 MUX2X1_254 ( .A(_1874_), .B(_1841_), .S(_1853__bF_buf2), .Y(_78__21_) );
INVX1 INVX1_1120 ( .A(_10732__22_), .Y(_1875_) );
MUX2X1 MUX2X1_255 ( .A(_1875_), .B(_1842_), .S(_1853__bF_buf1), .Y(_78__22_) );
INVX1 INVX1_1121 ( .A(_10732__23_), .Y(_1876_) );
MUX2X1 MUX2X1_256 ( .A(_1876_), .B(_1843_), .S(_1853__bF_buf0), .Y(_78__23_) );
INVX1 INVX1_1122 ( .A(_10732__24_), .Y(_1877_) );
NOR2X1 NOR2X1_1176 ( .A(_1853__bF_buf5), .B(_10728__24_), .Y(_1878_) );
AOI21X1 AOI21X1_874 ( .A(_1877_), .B(_1853__bF_buf4), .C(_1878_), .Y(_78__24_) );
INVX1 INVX1_1123 ( .A(_10732__25_), .Y(_1879_) );
NOR2X1 NOR2X1_1177 ( .A(_1853__bF_buf3), .B(_10728__25_), .Y(_1880_) );
AOI21X1 AOI21X1_875 ( .A(_1879_), .B(_1853__bF_buf2), .C(_1880_), .Y(_78__25_) );
INVX1 INVX1_1124 ( .A(_10732__26_), .Y(_1881_) );
NOR2X1 NOR2X1_1178 ( .A(_1853__bF_buf1), .B(_10728__26_), .Y(_1882_) );
AOI21X1 AOI21X1_876 ( .A(_1881_), .B(_1853__bF_buf0), .C(_1882_), .Y(_78__26_) );
INVX1 INVX1_1125 ( .A(_10732__27_), .Y(_1883_) );
NOR2X1 NOR2X1_1179 ( .A(_1853__bF_buf5), .B(_10728__27_), .Y(_1884_) );
AOI21X1 AOI21X1_877 ( .A(_1883_), .B(_1853__bF_buf4), .C(_1884_), .Y(_78__27_) );
INVX1 INVX1_1126 ( .A(_10732__28_), .Y(_1885_) );
NOR2X1 NOR2X1_1180 ( .A(_10728__28_), .B(_1853__bF_buf3), .Y(_1886_) );
AOI21X1 AOI21X1_878 ( .A(_1885_), .B(_1853__bF_buf2), .C(_1886_), .Y(_78__28_) );
INVX1 INVX1_1127 ( .A(_10732__29_), .Y(_1887_) );
NOR2X1 NOR2X1_1181 ( .A(_10728__29_), .B(_1853__bF_buf1), .Y(_1888_) );
AOI21X1 AOI21X1_879 ( .A(_1887_), .B(_1853__bF_buf0), .C(_1888_), .Y(_78__29_) );
INVX1 INVX1_1128 ( .A(_10732__30_), .Y(_1889_) );
NOR2X1 NOR2X1_1182 ( .A(_10728__30_), .B(_1853__bF_buf5), .Y(_1890_) );
AOI21X1 AOI21X1_880 ( .A(_1889_), .B(_1853__bF_buf4), .C(_1890_), .Y(_78__30_) );
INVX1 INVX1_1129 ( .A(_10732__31_), .Y(_1891_) );
NOR2X1 NOR2X1_1183 ( .A(_1853__bF_buf3), .B(_10728__31_), .Y(_1892_) );
AOI21X1 AOI21X1_881 ( .A(_1891_), .B(_1853__bF_buf2), .C(_1892_), .Y(_78__31_) );
OAI21X1 OAI21X1_2616 ( .A(_4937_), .B(_10103__bF_buf2), .C(_10130_), .Y(_1893_) );
OAI21X1 OAI21X1_2617 ( .A(mem_do_prefetch_bF_buf5), .B(mem_do_rinst_bF_buf4), .C(_1893_), .Y(_1894_) );
OAI21X1 OAI21X1_2618 ( .A(_5148_), .B(_4621__bF_buf2), .C(_1894_), .Y(_10726__2_) );
OAI21X1 OAI21X1_2619 ( .A(_4945_), .B(_10103__bF_buf1), .C(_10147_), .Y(_1895_) );
OAI21X1 OAI21X1_2620 ( .A(mem_do_prefetch_bF_buf4), .B(mem_do_rinst_bF_buf3), .C(_1895_), .Y(_1896_) );
OAI21X1 OAI21X1_2621 ( .A(_5130_), .B(_4621__bF_buf1), .C(_1896_), .Y(_10726__3_) );
OAI21X1 OAI21X1_2622 ( .A(_4952_), .B(_10103__bF_buf0), .C(_10165_), .Y(_1897_) );
OAI21X1 OAI21X1_2623 ( .A(mem_do_prefetch_bF_buf3), .B(mem_do_rinst_bF_buf2), .C(_1897_), .Y(_1898_) );
OAI21X1 OAI21X1_2624 ( .A(_5180_), .B(_4621__bF_buf0), .C(_1898_), .Y(_10726__4_) );
INVX1 INVX1_1130 ( .A(reg_out_5_), .Y(_1899_) );
OAI21X1 OAI21X1_2625 ( .A(_1899_), .B(_10103__bF_buf6), .C(_10191_), .Y(_1900_) );
OAI21X1 OAI21X1_2626 ( .A(mem_do_prefetch_bF_buf2), .B(mem_do_rinst_bF_buf1), .C(_1900_), .Y(_1901_) );
OAI21X1 OAI21X1_2627 ( .A(_5179_), .B(_4621__bF_buf4), .C(_1901_), .Y(_10726__5_) );
INVX1 INVX1_1131 ( .A(reg_out_6_), .Y(_1902_) );
OAI21X1 OAI21X1_2628 ( .A(_1902_), .B(_10103__bF_buf5), .C(_10205_), .Y(_1903_) );
OAI21X1 OAI21X1_2629 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf0), .C(_1903_), .Y(_1904_) );
OAI21X1 OAI21X1_2630 ( .A(_5174_), .B(_4621__bF_buf3), .C(_1904_), .Y(_10726__6_) );
INVX1 INVX1_1132 ( .A(reg_out_7_), .Y(_1905_) );
OAI21X1 OAI21X1_2631 ( .A(_1905_), .B(_10103__bF_buf4), .C(_10226_), .Y(_1906_) );
OAI21X1 OAI21X1_2632 ( .A(mem_do_prefetch_bF_buf0), .B(mem_do_rinst_bF_buf4), .C(_1906_), .Y(_1907_) );
OAI21X1 OAI21X1_2633 ( .A(_5173_), .B(_4621__bF_buf2), .C(_1907_), .Y(_10726__7_) );
INVX1 INVX1_1133 ( .A(reg_out_8_), .Y(_1908_) );
OAI21X1 OAI21X1_2634 ( .A(_1908_), .B(_10103__bF_buf3), .C(_10240_), .Y(_1909_) );
OAI21X1 OAI21X1_2635 ( .A(mem_do_prefetch_bF_buf5), .B(mem_do_rinst_bF_buf3), .C(_1909_), .Y(_1910_) );
OAI21X1 OAI21X1_2636 ( .A(_5187_), .B(_4621__bF_buf1), .C(_1910_), .Y(_10726__8_) );
OAI21X1 OAI21X1_2637 ( .A(_4693_), .B(_10103__bF_buf2), .C(_10271_), .Y(_1911_) );
OAI21X1 OAI21X1_2638 ( .A(mem_do_prefetch_bF_buf4), .B(mem_do_rinst_bF_buf2), .C(_1911_), .Y(_1912_) );
OAI21X1 OAI21X1_2639 ( .A(_5107_), .B(_4621__bF_buf0), .C(_1912_), .Y(_10726__9_) );
INVX1 INVX1_1134 ( .A(reg_out_10_), .Y(_1913_) );
OAI21X1 OAI21X1_2640 ( .A(_1913_), .B(_10103__bF_buf1), .C(_10284_), .Y(_1914_) );
OAI21X1 OAI21X1_2641 ( .A(mem_do_prefetch_bF_buf3), .B(mem_do_rinst_bF_buf1), .C(_1914_), .Y(_1915_) );
OAI21X1 OAI21X1_2642 ( .A(_5121_), .B(_4621__bF_buf4), .C(_1915_), .Y(_10726__10_) );
INVX1 INVX1_1135 ( .A(reg_out_11_), .Y(_1916_) );
OAI21X1 OAI21X1_2643 ( .A(_1916_), .B(_10103__bF_buf0), .C(_10314_), .Y(_1917_) );
OAI21X1 OAI21X1_2644 ( .A(mem_do_prefetch_bF_buf2), .B(mem_do_rinst_bF_buf0), .C(_1917_), .Y(_1918_) );
OAI21X1 OAI21X1_2645 ( .A(_5117_), .B(_4621__bF_buf3), .C(_1918_), .Y(_10726__11_) );
INVX1 INVX1_1136 ( .A(reg_out_12_), .Y(_1919_) );
OAI21X1 OAI21X1_2646 ( .A(_1919_), .B(_10103__bF_buf6), .C(_10330_), .Y(_1920_) );
OAI21X1 OAI21X1_2647 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf4), .C(_1920_), .Y(_1921_) );
OAI21X1 OAI21X1_2648 ( .A(_5197_), .B(_4621__bF_buf2), .C(_1921_), .Y(_10726__12_) );
OAI21X1 OAI21X1_2649 ( .A(_4724_), .B(_10103__bF_buf5), .C(_10364_), .Y(_1922_) );
OAI21X1 OAI21X1_2650 ( .A(mem_do_prefetch_bF_buf0), .B(mem_do_rinst_bF_buf3), .C(_1922_), .Y(_1923_) );
OAI21X1 OAI21X1_2651 ( .A(_5196_), .B(_4621__bF_buf1), .C(_1923_), .Y(_10726__13_) );
AOI21X1 AOI21X1_882 ( .A(reg_out_14_), .B(_10118__bF_buf0), .C(_10405_), .Y(_1924_) );
OAI21X1 OAI21X1_2652 ( .A(mem_do_prefetch_bF_buf5), .B(mem_do_rinst_bF_buf2), .C(_1924_), .Y(_1925_) );
OAI21X1 OAI21X1_2653 ( .A(_10734__14_), .B(_4621__bF_buf0), .C(_1925_), .Y(_1926_) );
INVX1 INVX1_1137 ( .A(_1926_), .Y(_10726__14_) );
INVX1 INVX1_1138 ( .A(reg_out_15_), .Y(_1927_) );
OAI21X1 OAI21X1_2654 ( .A(_1927_), .B(_10103__bF_buf4), .C(_10398_), .Y(_1928_) );
OAI21X1 OAI21X1_2655 ( .A(mem_do_prefetch_bF_buf4), .B(mem_do_rinst_bF_buf1), .C(_1928_), .Y(_1929_) );
OAI21X1 OAI21X1_2656 ( .A(_5087_), .B(_4621__bF_buf4), .C(_1929_), .Y(_10726__15_) );
OAI21X1 OAI21X1_2657 ( .A(_4749_), .B(_10103__bF_buf3), .C(_10429_), .Y(_1930_) );
OAI21X1 OAI21X1_2658 ( .A(mem_do_prefetch_bF_buf3), .B(mem_do_rinst_bF_buf0), .C(_1930_), .Y(_1931_) );
OAI21X1 OAI21X1_2659 ( .A(_5051_), .B(_4621__bF_buf3), .C(_1931_), .Y(_10726__16_) );
OAI21X1 OAI21X1_2660 ( .A(_4757_), .B(_10103__bF_buf2), .C(_10450_), .Y(_1932_) );
OAI21X1 OAI21X1_2661 ( .A(mem_do_prefetch_bF_buf2), .B(mem_do_rinst_bF_buf4), .C(_1932_), .Y(_1933_) );
OAI21X1 OAI21X1_2662 ( .A(_5057_), .B(_4621__bF_buf2), .C(_1933_), .Y(_10726__17_) );
OAI21X1 OAI21X1_2663 ( .A(_4765_), .B(_10103__bF_buf1), .C(_10472_), .Y(_1934_) );
OAI21X1 OAI21X1_2664 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf3), .C(_1934_), .Y(_1935_) );
OAI21X1 OAI21X1_2665 ( .A(_5045_), .B(_4621__bF_buf1), .C(_1935_), .Y(_10726__18_) );
INVX1 INVX1_1139 ( .A(_10491_), .Y(_1936_) );
OAI21X1 OAI21X1_2666 ( .A(_4785_), .B(_10103__bF_buf0), .C(_1936_), .Y(_1937_) );
OAI21X1 OAI21X1_2667 ( .A(mem_do_prefetch_bF_buf0), .B(mem_do_rinst_bF_buf2), .C(_1937_), .Y(_1938_) );
OAI21X1 OAI21X1_2668 ( .A(_5040_), .B(_4621__bF_buf0), .C(_1938_), .Y(_10726__19_) );
OAI21X1 OAI21X1_2669 ( .A(_10109__bF_buf3), .B(_4639__bF_buf0), .C(reg_next_pc_20_), .Y(_1939_) );
OAI21X1 OAI21X1_2670 ( .A(_4795_), .B(_10103__bF_buf6), .C(_1939_), .Y(_1940_) );
OAI21X1 OAI21X1_2671 ( .A(mem_do_prefetch_bF_buf5), .B(mem_do_rinst_bF_buf1), .C(_1940_), .Y(_1941_) );
OAI21X1 OAI21X1_2672 ( .A(_5218_), .B(_4621__bF_buf4), .C(_1941_), .Y(_10726__20_) );
OAI21X1 OAI21X1_2673 ( .A(_4808_), .B(_10103__bF_buf5), .C(_10542_), .Y(_1942_) );
OAI21X1 OAI21X1_2674 ( .A(mem_do_prefetch_bF_buf4), .B(mem_do_rinst_bF_buf0), .C(_1942_), .Y(_1943_) );
OAI21X1 OAI21X1_2675 ( .A(_5217_), .B(_4621__bF_buf3), .C(_1943_), .Y(_10726__21_) );
OAI21X1 OAI21X1_2676 ( .A(_10109__bF_buf2), .B(_4639__bF_buf4), .C(reg_next_pc_22_), .Y(_1944_) );
OAI21X1 OAI21X1_2677 ( .A(_4818_), .B(_10103__bF_buf4), .C(_1944_), .Y(_1945_) );
OAI21X1 OAI21X1_2678 ( .A(mem_do_prefetch_bF_buf3), .B(mem_do_rinst_bF_buf4), .C(_1945_), .Y(_1946_) );
OAI21X1 OAI21X1_2679 ( .A(_9021_), .B(_4621__bF_buf2), .C(_1946_), .Y(_10726__22_) );
OAI21X1 OAI21X1_2680 ( .A(_4828_), .B(_10103__bF_buf3), .C(_10586_), .Y(_1947_) );
OAI21X1 OAI21X1_2681 ( .A(mem_do_prefetch_bF_buf2), .B(mem_do_rinst_bF_buf3), .C(_1947_), .Y(_1948_) );
OAI21X1 OAI21X1_2682 ( .A(_9091_), .B(_4621__bF_buf1), .C(_1948_), .Y(_10726__23_) );
OAI21X1 OAI21X1_2683 ( .A(_4835_), .B(_10103__bF_buf2), .C(_10596_), .Y(_1949_) );
OAI21X1 OAI21X1_2684 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf2), .C(_1949_), .Y(_1950_) );
OAI21X1 OAI21X1_2685 ( .A(_5032_), .B(_4621__bF_buf0), .C(_1950_), .Y(_10726__24_) );
OAI21X1 OAI21X1_2686 ( .A(_4847_), .B(_10103__bF_buf1), .C(_10626_), .Y(_1951_) );
OAI21X1 OAI21X1_2687 ( .A(mem_do_prefetch_bF_buf0), .B(mem_do_rinst_bF_buf1), .C(_1951_), .Y(_1952_) );
OAI21X1 OAI21X1_2688 ( .A(_5027_), .B(_4621__bF_buf4), .C(_1952_), .Y(_10726__25_) );
OAI21X1 OAI21X1_2689 ( .A(_4856_), .B(_10103__bF_buf0), .C(_10644_), .Y(_1953_) );
OAI21X1 OAI21X1_2690 ( .A(mem_do_prefetch_bF_buf5), .B(mem_do_rinst_bF_buf0), .C(_1953_), .Y(_1954_) );
OAI21X1 OAI21X1_2691 ( .A(_5021_), .B(_4621__bF_buf3), .C(_1954_), .Y(_10726__26_) );
OAI21X1 OAI21X1_2692 ( .A(_4866_), .B(_10103__bF_buf6), .C(_10671_), .Y(_1955_) );
OAI21X1 OAI21X1_2693 ( .A(mem_do_prefetch_bF_buf4), .B(mem_do_rinst_bF_buf4), .C(_1955_), .Y(_1956_) );
OAI21X1 OAI21X1_2694 ( .A(_5016_), .B(_4621__bF_buf2), .C(_1956_), .Y(_10726__27_) );
OAI21X1 OAI21X1_2695 ( .A(_4873_), .B(_10103__bF_buf5), .C(_10686_), .Y(_1957_) );
OAI21X1 OAI21X1_2696 ( .A(mem_do_prefetch_bF_buf3), .B(mem_do_rinst_bF_buf3), .C(_1957_), .Y(_1958_) );
OAI21X1 OAI21X1_2697 ( .A(_5004_), .B(_4621__bF_buf1), .C(_1958_), .Y(_10726__28_) );
OAI21X1 OAI21X1_2698 ( .A(_4886_), .B(_10103__bF_buf4), .C(_10711_), .Y(_1959_) );
OAI21X1 OAI21X1_2699 ( .A(mem_do_prefetch_bF_buf2), .B(mem_do_rinst_bF_buf2), .C(_1959_), .Y(_1960_) );
OAI21X1 OAI21X1_2700 ( .A(_5009_), .B(_4621__bF_buf0), .C(_1960_), .Y(_10726__29_) );
OAI21X1 OAI21X1_2701 ( .A(_4895_), .B(_10103__bF_buf3), .C(_1128_), .Y(_1961_) );
OAI21X1 OAI21X1_2702 ( .A(mem_do_prefetch_bF_buf1), .B(mem_do_rinst_bF_buf1), .C(_1961_), .Y(_1962_) );
OAI21X1 OAI21X1_2703 ( .A(_4998_), .B(_4621__bF_buf4), .C(_1962_), .Y(_10726__30_) );
OAI21X1 OAI21X1_2704 ( .A(_4903_), .B(_10103__bF_buf2), .C(_1170_), .Y(_1963_) );
OAI21X1 OAI21X1_2705 ( .A(mem_do_prefetch_bF_buf0), .B(mem_do_rinst_bF_buf0), .C(_1963_), .Y(_1964_) );
OAI21X1 OAI21X1_2706 ( .A(_4991_), .B(_4621__bF_buf3), .C(_1964_), .Y(_10726__31_) );
INVX1 INVX1_1140 ( .A(_10724__0_), .Y(_1965_) );
INVX1 INVX1_1141 ( .A(_1782_), .Y(_1966_) );
NOR2X1 NOR2X1_1184 ( .A(_1966_), .B(_1802_), .Y(_1967_) );
NOR2X1 NOR2X1_1185 ( .A(_1965_), .B(_1967__bF_buf6), .Y(_70__0_) );
INVX1 INVX1_1142 ( .A(_10724__1_), .Y(_1968_) );
NOR2X1 NOR2X1_1186 ( .A(_1968_), .B(_1967__bF_buf5), .Y(_70__1_) );
INVX1 INVX1_1143 ( .A(_10726__2_), .Y(_1969_) );
NOR2X1 NOR2X1_1187 ( .A(_10724__2_), .B(_1967__bF_buf4), .Y(_1970_) );
AOI21X1 AOI21X1_883 ( .A(_1967__bF_buf3), .B(_1969_), .C(_1970_), .Y(_70__2_) );
INVX1 INVX1_1144 ( .A(_10726__3_), .Y(_1971_) );
NOR2X1 NOR2X1_1188 ( .A(_10724__3_), .B(_1967__bF_buf2), .Y(_1972_) );
AOI21X1 AOI21X1_884 ( .A(_1967__bF_buf1), .B(_1971_), .C(_1972_), .Y(_70__3_) );
INVX1 INVX1_1145 ( .A(_10726__4_), .Y(_1973_) );
NOR2X1 NOR2X1_1189 ( .A(_10724__4_), .B(_1967__bF_buf0), .Y(_1974_) );
AOI21X1 AOI21X1_885 ( .A(_1967__bF_buf6), .B(_1973_), .C(_1974_), .Y(_70__4_) );
INVX1 INVX1_1146 ( .A(_10726__5_), .Y(_1975_) );
NOR2X1 NOR2X1_1190 ( .A(_10724__5_), .B(_1967__bF_buf5), .Y(_1976_) );
AOI21X1 AOI21X1_886 ( .A(_1967__bF_buf4), .B(_1975_), .C(_1976_), .Y(_70__5_) );
INVX1 INVX1_1147 ( .A(_10726__6_), .Y(_1977_) );
NOR2X1 NOR2X1_1191 ( .A(_10724__6_), .B(_1967__bF_buf3), .Y(_1978_) );
AOI21X1 AOI21X1_887 ( .A(_1967__bF_buf2), .B(_1977_), .C(_1978_), .Y(_70__6_) );
INVX1 INVX1_1148 ( .A(_10726__7_), .Y(_1979_) );
NOR2X1 NOR2X1_1192 ( .A(_10724__7_), .B(_1967__bF_buf1), .Y(_1980_) );
AOI21X1 AOI21X1_888 ( .A(_1967__bF_buf0), .B(_1979_), .C(_1980_), .Y(_70__7_) );
INVX1 INVX1_1149 ( .A(_10726__8_), .Y(_1981_) );
NOR2X1 NOR2X1_1193 ( .A(_10724__8_), .B(_1967__bF_buf6), .Y(_1982_) );
AOI21X1 AOI21X1_889 ( .A(_1967__bF_buf5), .B(_1981_), .C(_1982_), .Y(_70__8_) );
INVX1 INVX1_1150 ( .A(_10726__9_), .Y(_1983_) );
NOR2X1 NOR2X1_1194 ( .A(_10724__9_), .B(_1967__bF_buf4), .Y(_1984_) );
AOI21X1 AOI21X1_890 ( .A(_1967__bF_buf3), .B(_1983_), .C(_1984_), .Y(_70__9_) );
INVX1 INVX1_1151 ( .A(_10726__10_), .Y(_1985_) );
NOR2X1 NOR2X1_1195 ( .A(_10724__10_), .B(_1967__bF_buf2), .Y(_1986_) );
AOI21X1 AOI21X1_891 ( .A(_1967__bF_buf1), .B(_1985_), .C(_1986_), .Y(_70__10_) );
INVX1 INVX1_1152 ( .A(_10726__11_), .Y(_1987_) );
NOR2X1 NOR2X1_1196 ( .A(_10724__11_), .B(_1967__bF_buf0), .Y(_1988_) );
AOI21X1 AOI21X1_892 ( .A(_1967__bF_buf6), .B(_1987_), .C(_1988_), .Y(_70__11_) );
INVX1 INVX1_1153 ( .A(_10726__12_), .Y(_1989_) );
NOR2X1 NOR2X1_1197 ( .A(_10724__12_), .B(_1967__bF_buf5), .Y(_1990_) );
AOI21X1 AOI21X1_893 ( .A(_1967__bF_buf4), .B(_1989_), .C(_1990_), .Y(_70__12_) );
INVX1 INVX1_1154 ( .A(_10726__13_), .Y(_1991_) );
NOR2X1 NOR2X1_1198 ( .A(_10724__13_), .B(_1967__bF_buf3), .Y(_1992_) );
AOI21X1 AOI21X1_894 ( .A(_1967__bF_buf2), .B(_1991_), .C(_1992_), .Y(_70__13_) );
NOR2X1 NOR2X1_1199 ( .A(_10724__14_), .B(_1967__bF_buf1), .Y(_1993_) );
AOI21X1 AOI21X1_895 ( .A(_1967__bF_buf0), .B(_1926_), .C(_1993_), .Y(_70__14_) );
INVX1 INVX1_1155 ( .A(_10726__15_), .Y(_1994_) );
NOR2X1 NOR2X1_1200 ( .A(_10724__15_), .B(_1967__bF_buf6), .Y(_1995_) );
AOI21X1 AOI21X1_896 ( .A(_1967__bF_buf5), .B(_1994_), .C(_1995_), .Y(_70__15_) );
INVX1 INVX1_1156 ( .A(_10726__16_), .Y(_1996_) );
NOR2X1 NOR2X1_1201 ( .A(_10724__16_), .B(_1967__bF_buf4), .Y(_1997_) );
AOI21X1 AOI21X1_897 ( .A(_1967__bF_buf3), .B(_1996_), .C(_1997_), .Y(_70__16_) );
INVX1 INVX1_1157 ( .A(_10726__17_), .Y(_1998_) );
NOR2X1 NOR2X1_1202 ( .A(_10724__17_), .B(_1967__bF_buf2), .Y(_1999_) );
AOI21X1 AOI21X1_898 ( .A(_1967__bF_buf1), .B(_1998_), .C(_1999_), .Y(_70__17_) );
INVX1 INVX1_1158 ( .A(_10726__18_), .Y(_2000_) );
NOR2X1 NOR2X1_1203 ( .A(_10724__18_), .B(_1967__bF_buf0), .Y(_2001_) );
AOI21X1 AOI21X1_899 ( .A(_1967__bF_buf6), .B(_2000_), .C(_2001_), .Y(_70__18_) );
INVX1 INVX1_1159 ( .A(_10726__19_), .Y(_2002_) );
NOR2X1 NOR2X1_1204 ( .A(_10724__19_), .B(_1967__bF_buf5), .Y(_2003_) );
AOI21X1 AOI21X1_900 ( .A(_1967__bF_buf4), .B(_2002_), .C(_2003_), .Y(_70__19_) );
INVX1 INVX1_1160 ( .A(_10726__20_), .Y(_2004_) );
NOR2X1 NOR2X1_1205 ( .A(_10724__20_), .B(_1967__bF_buf3), .Y(_2005_) );
AOI21X1 AOI21X1_901 ( .A(_1967__bF_buf2), .B(_2004_), .C(_2005_), .Y(_70__20_) );
INVX1 INVX1_1161 ( .A(_10726__21_), .Y(_2006_) );
NOR2X1 NOR2X1_1206 ( .A(_10724__21_), .B(_1967__bF_buf1), .Y(_2007_) );
AOI21X1 AOI21X1_902 ( .A(_1967__bF_buf0), .B(_2006_), .C(_2007_), .Y(_70__21_) );
INVX1 INVX1_1162 ( .A(_10726__22_), .Y(_2008_) );
NOR2X1 NOR2X1_1207 ( .A(_10724__22_), .B(_1967__bF_buf6), .Y(_2009_) );
AOI21X1 AOI21X1_903 ( .A(_1967__bF_buf5), .B(_2008_), .C(_2009_), .Y(_70__22_) );
INVX1 INVX1_1163 ( .A(_10726__23_), .Y(_2010_) );
NOR2X1 NOR2X1_1208 ( .A(_10724__23_), .B(_1967__bF_buf4), .Y(_2011_) );
AOI21X1 AOI21X1_904 ( .A(_1967__bF_buf3), .B(_2010_), .C(_2011_), .Y(_70__23_) );
INVX1 INVX1_1164 ( .A(_10726__24_), .Y(_2012_) );
NOR2X1 NOR2X1_1209 ( .A(_10724__24_), .B(_1967__bF_buf2), .Y(_2013_) );
AOI21X1 AOI21X1_905 ( .A(_1967__bF_buf1), .B(_2012_), .C(_2013_), .Y(_70__24_) );
INVX1 INVX1_1165 ( .A(_10726__25_), .Y(_2014_) );
NOR2X1 NOR2X1_1210 ( .A(_10724__25_), .B(_1967__bF_buf0), .Y(_2015_) );
AOI21X1 AOI21X1_906 ( .A(_1967__bF_buf6), .B(_2014_), .C(_2015_), .Y(_70__25_) );
INVX1 INVX1_1166 ( .A(_10726__26_), .Y(_2016_) );
NOR2X1 NOR2X1_1211 ( .A(_10724__26_), .B(_1967__bF_buf5), .Y(_2017_) );
AOI21X1 AOI21X1_907 ( .A(_1967__bF_buf4), .B(_2016_), .C(_2017_), .Y(_70__26_) );
INVX1 INVX1_1167 ( .A(_10726__27_), .Y(_2018_) );
NOR2X1 NOR2X1_1212 ( .A(_10724__27_), .B(_1967__bF_buf3), .Y(_2019_) );
AOI21X1 AOI21X1_908 ( .A(_1967__bF_buf2), .B(_2018_), .C(_2019_), .Y(_70__27_) );
INVX1 INVX1_1168 ( .A(_10726__28_), .Y(_2020_) );
NOR2X1 NOR2X1_1213 ( .A(_10724__28_), .B(_1967__bF_buf1), .Y(_2021_) );
AOI21X1 AOI21X1_909 ( .A(_1967__bF_buf0), .B(_2020_), .C(_2021_), .Y(_70__28_) );
INVX1 INVX1_1169 ( .A(_10726__29_), .Y(_2022_) );
NOR2X1 NOR2X1_1214 ( .A(_10724__29_), .B(_1967__bF_buf6), .Y(_2023_) );
AOI21X1 AOI21X1_910 ( .A(_1967__bF_buf5), .B(_2022_), .C(_2023_), .Y(_70__29_) );
INVX1 INVX1_1170 ( .A(_10726__30_), .Y(_2024_) );
NOR2X1 NOR2X1_1215 ( .A(_10724__30_), .B(_1967__bF_buf4), .Y(_2025_) );
AOI21X1 AOI21X1_911 ( .A(_1967__bF_buf3), .B(_2024_), .C(_2025_), .Y(_70__30_) );
INVX1 INVX1_1171 ( .A(_10726__31_), .Y(_2026_) );
NOR2X1 NOR2X1_1216 ( .A(_10724__31_), .B(_1967__bF_buf2), .Y(_2027_) );
AOI21X1 AOI21X1_912 ( .A(_1967__bF_buf1), .B(_2026_), .C(_2027_), .Y(_70__31_) );
AOI22X1 AOI22X1_128 ( .A(_4427_), .B(_10725_), .C(_4621__bF_buf2), .D(_1782_), .Y(_2028_) );
OAI21X1 OAI21X1_2707 ( .A(_1966_), .B(_4619_), .C(_10725_), .Y(_2029_) );
OAI21X1 OAI21X1_2708 ( .A(_1784_), .B(_2028_), .C(_2029_), .Y(_75_) );
OAI21X1 OAI21X1_2709 ( .A(_4619_), .B(_10736_), .C(resetn_bF_buf1), .Y(_2030_) );
OAI21X1 OAI21X1_2710 ( .A(_4434_), .B(_4438_), .C(_1782_), .Y(_2031_) );
OAI21X1 OAI21X1_2711 ( .A(_2030_), .B(mem_ready), .C(_2031_), .Y(_2032_) );
NAND2X1 NAND2X1_890 ( .A(_10731_), .B(_2032_), .Y(_2033_) );
OAI21X1 OAI21X1_2712 ( .A(_1802_), .B(_1966_), .C(_2033_), .Y(_77_) );
NOR2X1 NOR2X1_1217 ( .A(_4633_), .B(_5743_), .Y(_2034_) );
NAND2X1 NAND2X1_891 ( .A(latched_rd_2_), .B(_2034_), .Y(_2035_) );
INVX1 INVX1_1172 ( .A(_2035__bF_buf8), .Y(_2036_) );
NAND2X1 NAND2X1_892 ( .A(_2036_), .B(_5745_), .Y(_2037_) );
OAI21X1 OAI21X1_2713 ( .A(_4917__bF_buf9), .B(_2035__bF_buf7), .C(cpuregs_31_[0]), .Y(_2038_) );
OAI21X1 OAI21X1_2714 ( .A(_2037__bF_buf4), .B(_4925__bF_buf2), .C(_2038_), .Y(_379_) );
OAI21X1 OAI21X1_2715 ( .A(_4917__bF_buf8), .B(_2035__bF_buf6), .C(cpuregs_31_[1]), .Y(_2039_) );
OAI21X1 OAI21X1_2716 ( .A(_2037__bF_buf3), .B(_4933__bF_buf2), .C(_2039_), .Y(_380_) );
OAI21X1 OAI21X1_2717 ( .A(_4917__bF_buf7), .B(_2035__bF_buf5), .C(cpuregs_31_[2]), .Y(_2040_) );
OAI21X1 OAI21X1_2718 ( .A(_2037__bF_buf2), .B(_4940__bF_buf2), .C(_2040_), .Y(_381_) );
OAI21X1 OAI21X1_2719 ( .A(_4917__bF_buf6), .B(_2035__bF_buf4), .C(cpuregs_31_[3]), .Y(_2041_) );
OAI21X1 OAI21X1_2720 ( .A(_2037__bF_buf1), .B(_4948__bF_buf2), .C(_2041_), .Y(_382_) );
OAI21X1 OAI21X1_2721 ( .A(_4917__bF_buf5), .B(_2035__bF_buf3), .C(cpuregs_31_[4]), .Y(_2042_) );
OAI21X1 OAI21X1_2722 ( .A(_2037__bF_buf0), .B(_4955__bF_buf2), .C(_2042_), .Y(_383_) );
OAI21X1 OAI21X1_2723 ( .A(_4917__bF_buf4), .B(_2035__bF_buf2), .C(cpuregs_31_[5]), .Y(_2043_) );
OAI21X1 OAI21X1_2724 ( .A(_2037__bF_buf4), .B(_4654__bF_buf1), .C(_2043_), .Y(_384_) );
OAI21X1 OAI21X1_2725 ( .A(_4917__bF_buf3), .B(_2035__bF_buf1), .C(cpuregs_31_[6]), .Y(_2044_) );
OAI21X1 OAI21X1_2726 ( .A(_4664__bF_buf1), .B(_2037__bF_buf3), .C(_2044_), .Y(_385_) );
OAI21X1 OAI21X1_2727 ( .A(_4917__bF_buf2), .B(_2035__bF_buf0), .C(cpuregs_31_[7]), .Y(_2045_) );
OAI21X1 OAI21X1_2728 ( .A(_4677__bF_buf1), .B(_2037__bF_buf2), .C(_2045_), .Y(_386_) );
OAI21X1 OAI21X1_2729 ( .A(_4917__bF_buf1), .B(_2035__bF_buf8), .C(cpuregs_31_[8]), .Y(_2046_) );
OAI21X1 OAI21X1_2730 ( .A(_4685__bF_buf1), .B(_2037__bF_buf1), .C(_2046_), .Y(_387_) );
OAI21X1 OAI21X1_2731 ( .A(_4917__bF_buf0), .B(_2035__bF_buf7), .C(cpuregs_31_[9]), .Y(_2047_) );
OAI21X1 OAI21X1_2732 ( .A(_4696__bF_buf1), .B(_2037__bF_buf0), .C(_2047_), .Y(_388_) );
OAI21X1 OAI21X1_2733 ( .A(_4917__bF_buf10), .B(_2035__bF_buf6), .C(cpuregs_31_[10]), .Y(_2048_) );
OAI21X1 OAI21X1_2734 ( .A(_4703__bF_buf1), .B(_2037__bF_buf4), .C(_2048_), .Y(_389_) );
OAI21X1 OAI21X1_2735 ( .A(_4917__bF_buf9), .B(_2035__bF_buf5), .C(cpuregs_31_[11]), .Y(_2049_) );
OAI21X1 OAI21X1_2736 ( .A(_4713__bF_buf1), .B(_2037__bF_buf3), .C(_2049_), .Y(_390_) );
OAI21X1 OAI21X1_2737 ( .A(_4917__bF_buf8), .B(_2035__bF_buf4), .C(cpuregs_31_[12]), .Y(_2050_) );
OAI21X1 OAI21X1_2738 ( .A(_4722__bF_buf1), .B(_2037__bF_buf2), .C(_2050_), .Y(_391_) );
OAI21X1 OAI21X1_2739 ( .A(_4917__bF_buf7), .B(_2035__bF_buf3), .C(cpuregs_31_[13]), .Y(_2051_) );
OAI21X1 OAI21X1_2740 ( .A(_4731__bF_buf1), .B(_2037__bF_buf1), .C(_2051_), .Y(_392_) );
OAI21X1 OAI21X1_2741 ( .A(_4917__bF_buf6), .B(_2035__bF_buf2), .C(cpuregs_31_[14]), .Y(_2052_) );
OAI21X1 OAI21X1_2742 ( .A(_4740__bF_buf1), .B(_2037__bF_buf0), .C(_2052_), .Y(_393_) );
OAI21X1 OAI21X1_2743 ( .A(_4917__bF_buf5), .B(_2035__bF_buf1), .C(cpuregs_31_[15]), .Y(_2053_) );
OAI21X1 OAI21X1_2744 ( .A(_4747__bF_buf1), .B(_2037__bF_buf4), .C(_2053_), .Y(_394_) );
OAI21X1 OAI21X1_2745 ( .A(_4917__bF_buf4), .B(_2035__bF_buf0), .C(cpuregs_31_[16]), .Y(_2054_) );
OAI21X1 OAI21X1_2746 ( .A(_4755__bF_buf1), .B(_2037__bF_buf3), .C(_2054_), .Y(_395_) );
OAI21X1 OAI21X1_2747 ( .A(_4917__bF_buf3), .B(_2035__bF_buf8), .C(cpuregs_31_[17]), .Y(_2055_) );
OAI21X1 OAI21X1_2748 ( .A(_4763__bF_buf1), .B(_2037__bF_buf2), .C(_2055_), .Y(_396_) );
OAI21X1 OAI21X1_2749 ( .A(_4917__bF_buf2), .B(_2035__bF_buf7), .C(cpuregs_31_[18]), .Y(_2056_) );
OAI21X1 OAI21X1_2750 ( .A(_4783__bF_buf1), .B(_2037__bF_buf1), .C(_2056_), .Y(_397_) );
OAI21X1 OAI21X1_2751 ( .A(_4917__bF_buf1), .B(_2035__bF_buf6), .C(cpuregs_31_[19]), .Y(_2057_) );
OAI21X1 OAI21X1_2752 ( .A(_4793__bF_buf1), .B(_2037__bF_buf0), .C(_2057_), .Y(_398_) );
OAI21X1 OAI21X1_2753 ( .A(_4917__bF_buf0), .B(_2035__bF_buf5), .C(cpuregs_31_[20]), .Y(_2058_) );
OAI21X1 OAI21X1_2754 ( .A(_4806__bF_buf1), .B(_2037__bF_buf4), .C(_2058_), .Y(_399_) );
OAI21X1 OAI21X1_2755 ( .A(_4917__bF_buf10), .B(_2035__bF_buf4), .C(cpuregs_31_[21]), .Y(_2059_) );
OAI21X1 OAI21X1_2756 ( .A(_4816__bF_buf1), .B(_2037__bF_buf3), .C(_2059_), .Y(_400_) );
OAI21X1 OAI21X1_2757 ( .A(_4917__bF_buf9), .B(_2035__bF_buf3), .C(cpuregs_31_[22]), .Y(_2060_) );
OAI21X1 OAI21X1_2758 ( .A(_4824__bF_buf1), .B(_2037__bF_buf2), .C(_2060_), .Y(_401_) );
OAI21X1 OAI21X1_2759 ( .A(_4917__bF_buf8), .B(_2035__bF_buf2), .C(cpuregs_31_[23]), .Y(_2061_) );
OAI21X1 OAI21X1_2760 ( .A(_4833__bF_buf1), .B(_2037__bF_buf1), .C(_2061_), .Y(_402_) );
OAI21X1 OAI21X1_2761 ( .A(_4917__bF_buf7), .B(_2035__bF_buf1), .C(cpuregs_31_[24]), .Y(_2062_) );
OAI21X1 OAI21X1_2762 ( .A(_4845__bF_buf1), .B(_2037__bF_buf0), .C(_2062_), .Y(_403_) );
OAI21X1 OAI21X1_2763 ( .A(_4917__bF_buf6), .B(_2035__bF_buf0), .C(cpuregs_31_[25]), .Y(_2063_) );
OAI21X1 OAI21X1_2764 ( .A(_4854__bF_buf1), .B(_2037__bF_buf4), .C(_2063_), .Y(_404_) );
OAI21X1 OAI21X1_2765 ( .A(_4917__bF_buf5), .B(_2035__bF_buf8), .C(cpuregs_31_[26]), .Y(_2064_) );
OAI21X1 OAI21X1_2766 ( .A(_4863__bF_buf1), .B(_2037__bF_buf3), .C(_2064_), .Y(_405_) );
OAI21X1 OAI21X1_2767 ( .A(_4917__bF_buf4), .B(_2035__bF_buf7), .C(cpuregs_31_[27]), .Y(_2065_) );
OAI21X1 OAI21X1_2768 ( .A(_4871__bF_buf1), .B(_2037__bF_buf2), .C(_2065_), .Y(_406_) );
OAI21X1 OAI21X1_2769 ( .A(_4917__bF_buf3), .B(_2035__bF_buf6), .C(cpuregs_31_[28]), .Y(_2066_) );
OAI21X1 OAI21X1_2770 ( .A(_4884__bF_buf1), .B(_2037__bF_buf1), .C(_2066_), .Y(_407_) );
OAI21X1 OAI21X1_2771 ( .A(_4917__bF_buf2), .B(_2035__bF_buf5), .C(cpuregs_31_[29]), .Y(_2067_) );
OAI21X1 OAI21X1_2772 ( .A(_4893__bF_buf1), .B(_2037__bF_buf0), .C(_2067_), .Y(_408_) );
OAI21X1 OAI21X1_2773 ( .A(_4917__bF_buf1), .B(_2035__bF_buf4), .C(cpuregs_31_[30]), .Y(_2068_) );
OAI21X1 OAI21X1_2774 ( .A(_4901__bF_buf1), .B(_2037__bF_buf4), .C(_2068_), .Y(_409_) );
OAI21X1 OAI21X1_2775 ( .A(_4917__bF_buf0), .B(_2035__bF_buf3), .C(cpuregs_31_[31]), .Y(_2069_) );
OAI21X1 OAI21X1_2776 ( .A(_4910__bF_buf1), .B(_2037__bF_buf3), .C(_2069_), .Y(_410_) );
NOR2X1 NOR2X1_1218 ( .A(_2035__bF_buf2), .B(_5281__bF_buf8), .Y(_2070_) );
INVX1 INVX1_1173 ( .A(_2070_), .Y(_2071_) );
OAI21X1 OAI21X1_2777 ( .A(_5281__bF_buf7), .B(_2035__bF_buf1), .C(cpuregs_30_[0]), .Y(_2072_) );
OAI21X1 OAI21X1_2778 ( .A(_2071__bF_buf4), .B(_4925__bF_buf1), .C(_2072_), .Y(_411_) );
OAI21X1 OAI21X1_2779 ( .A(_5281__bF_buf6), .B(_2035__bF_buf0), .C(cpuregs_30_[1]), .Y(_2073_) );
OAI21X1 OAI21X1_2780 ( .A(_2071__bF_buf3), .B(_4933__bF_buf1), .C(_2073_), .Y(_412_) );
OAI21X1 OAI21X1_2781 ( .A(_5281__bF_buf5), .B(_2035__bF_buf8), .C(cpuregs_30_[2]), .Y(_2074_) );
OAI21X1 OAI21X1_2782 ( .A(_2071__bF_buf2), .B(_4940__bF_buf1), .C(_2074_), .Y(_413_) );
OAI21X1 OAI21X1_2783 ( .A(_5281__bF_buf4), .B(_2035__bF_buf7), .C(cpuregs_30_[3]), .Y(_2075_) );
OAI21X1 OAI21X1_2784 ( .A(_2071__bF_buf1), .B(_4948__bF_buf1), .C(_2075_), .Y(_414_) );
OAI21X1 OAI21X1_2785 ( .A(_5281__bF_buf3), .B(_2035__bF_buf6), .C(cpuregs_30_[4]), .Y(_2076_) );
OAI21X1 OAI21X1_2786 ( .A(_2071__bF_buf0), .B(_4955__bF_buf1), .C(_2076_), .Y(_415_) );
OAI21X1 OAI21X1_2787 ( .A(_5281__bF_buf2), .B(_2035__bF_buf5), .C(cpuregs_30_[5]), .Y(_2077_) );
OAI21X1 OAI21X1_2788 ( .A(_2071__bF_buf4), .B(_4654__bF_buf0), .C(_2077_), .Y(_416_) );
OAI21X1 OAI21X1_2789 ( .A(_5281__bF_buf1), .B(_2035__bF_buf4), .C(cpuregs_30_[6]), .Y(_2078_) );
OAI21X1 OAI21X1_2790 ( .A(_4664__bF_buf0), .B(_2071__bF_buf3), .C(_2078_), .Y(_417_) );
OAI21X1 OAI21X1_2791 ( .A(_5281__bF_buf0), .B(_2035__bF_buf3), .C(cpuregs_30_[7]), .Y(_2079_) );
OAI21X1 OAI21X1_2792 ( .A(_4677__bF_buf0), .B(_2071__bF_buf2), .C(_2079_), .Y(_418_) );
OAI21X1 OAI21X1_2793 ( .A(_5281__bF_buf10), .B(_2035__bF_buf2), .C(cpuregs_30_[8]), .Y(_2080_) );
OAI21X1 OAI21X1_2794 ( .A(_4685__bF_buf0), .B(_2071__bF_buf1), .C(_2080_), .Y(_419_) );
OAI21X1 OAI21X1_2795 ( .A(_5281__bF_buf9), .B(_2035__bF_buf1), .C(cpuregs_30_[9]), .Y(_2081_) );
OAI21X1 OAI21X1_2796 ( .A(_4696__bF_buf0), .B(_2071__bF_buf0), .C(_2081_), .Y(_420_) );
OAI21X1 OAI21X1_2797 ( .A(_5281__bF_buf8), .B(_2035__bF_buf0), .C(cpuregs_30_[10]), .Y(_2082_) );
OAI21X1 OAI21X1_2798 ( .A(_4703__bF_buf0), .B(_2071__bF_buf4), .C(_2082_), .Y(_421_) );
OAI21X1 OAI21X1_2799 ( .A(_5281__bF_buf7), .B(_2035__bF_buf8), .C(cpuregs_30_[11]), .Y(_2083_) );
OAI21X1 OAI21X1_2800 ( .A(_4713__bF_buf0), .B(_2071__bF_buf3), .C(_2083_), .Y(_422_) );
OAI21X1 OAI21X1_2801 ( .A(_5281__bF_buf6), .B(_2035__bF_buf7), .C(cpuregs_30_[12]), .Y(_2084_) );
OAI21X1 OAI21X1_2802 ( .A(_4722__bF_buf0), .B(_2071__bF_buf2), .C(_2084_), .Y(_423_) );
OAI21X1 OAI21X1_2803 ( .A(_5281__bF_buf5), .B(_2035__bF_buf6), .C(cpuregs_30_[13]), .Y(_2085_) );
OAI21X1 OAI21X1_2804 ( .A(_4731__bF_buf0), .B(_2071__bF_buf1), .C(_2085_), .Y(_424_) );
OAI21X1 OAI21X1_2805 ( .A(_5281__bF_buf4), .B(_2035__bF_buf5), .C(cpuregs_30_[14]), .Y(_2086_) );
OAI21X1 OAI21X1_2806 ( .A(_4740__bF_buf0), .B(_2071__bF_buf0), .C(_2086_), .Y(_425_) );
OAI21X1 OAI21X1_2807 ( .A(_5281__bF_buf3), .B(_2035__bF_buf4), .C(cpuregs_30_[15]), .Y(_2087_) );
OAI21X1 OAI21X1_2808 ( .A(_4747__bF_buf0), .B(_2071__bF_buf4), .C(_2087_), .Y(_426_) );
OAI21X1 OAI21X1_2809 ( .A(_5281__bF_buf2), .B(_2035__bF_buf3), .C(cpuregs_30_[16]), .Y(_2088_) );
OAI21X1 OAI21X1_2810 ( .A(_4755__bF_buf0), .B(_2071__bF_buf3), .C(_2088_), .Y(_427_) );
OAI21X1 OAI21X1_2811 ( .A(_5281__bF_buf1), .B(_2035__bF_buf2), .C(cpuregs_30_[17]), .Y(_2089_) );
OAI21X1 OAI21X1_2812 ( .A(_4763__bF_buf0), .B(_2071__bF_buf2), .C(_2089_), .Y(_428_) );
OAI21X1 OAI21X1_2813 ( .A(_5281__bF_buf0), .B(_2035__bF_buf1), .C(cpuregs_30_[18]), .Y(_2090_) );
OAI21X1 OAI21X1_2814 ( .A(_4783__bF_buf0), .B(_2071__bF_buf1), .C(_2090_), .Y(_429_) );
OAI21X1 OAI21X1_2815 ( .A(_5281__bF_buf10), .B(_2035__bF_buf0), .C(cpuregs_30_[19]), .Y(_2091_) );
OAI21X1 OAI21X1_2816 ( .A(_4793__bF_buf0), .B(_2071__bF_buf0), .C(_2091_), .Y(_430_) );
OAI21X1 OAI21X1_2817 ( .A(_5281__bF_buf9), .B(_2035__bF_buf8), .C(cpuregs_30_[20]), .Y(_2092_) );
OAI21X1 OAI21X1_2818 ( .A(_4806__bF_buf0), .B(_2071__bF_buf4), .C(_2092_), .Y(_431_) );
OAI21X1 OAI21X1_2819 ( .A(_5281__bF_buf8), .B(_2035__bF_buf7), .C(cpuregs_30_[21]), .Y(_2093_) );
OAI21X1 OAI21X1_2820 ( .A(_4816__bF_buf0), .B(_2071__bF_buf3), .C(_2093_), .Y(_432_) );
OAI21X1 OAI21X1_2821 ( .A(_5281__bF_buf7), .B(_2035__bF_buf6), .C(cpuregs_30_[22]), .Y(_2094_) );
OAI21X1 OAI21X1_2822 ( .A(_4824__bF_buf0), .B(_2071__bF_buf2), .C(_2094_), .Y(_433_) );
OAI21X1 OAI21X1_2823 ( .A(_5281__bF_buf6), .B(_2035__bF_buf5), .C(cpuregs_30_[23]), .Y(_2095_) );
OAI21X1 OAI21X1_2824 ( .A(_4833__bF_buf0), .B(_2071__bF_buf1), .C(_2095_), .Y(_434_) );
OAI21X1 OAI21X1_2825 ( .A(_5281__bF_buf5), .B(_2035__bF_buf4), .C(cpuregs_30_[24]), .Y(_2096_) );
OAI21X1 OAI21X1_2826 ( .A(_4845__bF_buf0), .B(_2071__bF_buf0), .C(_2096_), .Y(_435_) );
OAI21X1 OAI21X1_2827 ( .A(_5281__bF_buf4), .B(_2035__bF_buf3), .C(cpuregs_30_[25]), .Y(_2097_) );
OAI21X1 OAI21X1_2828 ( .A(_4854__bF_buf0), .B(_2071__bF_buf4), .C(_2097_), .Y(_436_) );
OAI21X1 OAI21X1_2829 ( .A(_5281__bF_buf3), .B(_2035__bF_buf2), .C(cpuregs_30_[26]), .Y(_2098_) );
OAI21X1 OAI21X1_2830 ( .A(_4863__bF_buf0), .B(_2071__bF_buf3), .C(_2098_), .Y(_437_) );
OAI21X1 OAI21X1_2831 ( .A(_5281__bF_buf2), .B(_2035__bF_buf1), .C(cpuregs_30_[27]), .Y(_2099_) );
OAI21X1 OAI21X1_2832 ( .A(_4871__bF_buf0), .B(_2071__bF_buf2), .C(_2099_), .Y(_438_) );
OAI21X1 OAI21X1_2833 ( .A(_5281__bF_buf1), .B(_2035__bF_buf0), .C(cpuregs_30_[28]), .Y(_2100_) );
OAI21X1 OAI21X1_2834 ( .A(_4884__bF_buf0), .B(_2071__bF_buf1), .C(_2100_), .Y(_439_) );
OAI21X1 OAI21X1_2835 ( .A(_5281__bF_buf0), .B(_2035__bF_buf8), .C(cpuregs_30_[29]), .Y(_2101_) );
OAI21X1 OAI21X1_2836 ( .A(_4893__bF_buf0), .B(_2071__bF_buf0), .C(_2101_), .Y(_440_) );
OAI21X1 OAI21X1_2837 ( .A(_5281__bF_buf10), .B(_2035__bF_buf7), .C(cpuregs_30_[30]), .Y(_2102_) );
OAI21X1 OAI21X1_2838 ( .A(_4901__bF_buf0), .B(_2071__bF_buf4), .C(_2102_), .Y(_441_) );
OAI21X1 OAI21X1_2839 ( .A(_5281__bF_buf9), .B(_2035__bF_buf6), .C(cpuregs_30_[31]), .Y(_2103_) );
OAI21X1 OAI21X1_2840 ( .A(_4910__bF_buf0), .B(_2071__bF_buf3), .C(_2103_), .Y(_442_) );
NAND2X1 NAND2X1_893 ( .A(_2036_), .B(_5313_), .Y(_2104_) );
NAND2X1 NAND2X1_894 ( .A(cpuregs_29_[0]), .B(_2104__bF_buf7), .Y(_2105_) );
OAI21X1 OAI21X1_2841 ( .A(_4925__bF_buf0), .B(_2104__bF_buf6), .C(_2105_), .Y(_443_) );
NAND2X1 NAND2X1_895 ( .A(cpuregs_29_[1]), .B(_2104__bF_buf5), .Y(_2106_) );
OAI21X1 OAI21X1_2842 ( .A(_4933__bF_buf0), .B(_2104__bF_buf4), .C(_2106_), .Y(_444_) );
NAND2X1 NAND2X1_896 ( .A(cpuregs_29_[2]), .B(_2104__bF_buf3), .Y(_2107_) );
OAI21X1 OAI21X1_2843 ( .A(_4940__bF_buf0), .B(_2104__bF_buf2), .C(_2107_), .Y(_445_) );
NAND2X1 NAND2X1_897 ( .A(cpuregs_29_[3]), .B(_2104__bF_buf1), .Y(_2108_) );
OAI21X1 OAI21X1_2844 ( .A(_4948__bF_buf0), .B(_2104__bF_buf0), .C(_2108_), .Y(_446_) );
NAND2X1 NAND2X1_898 ( .A(cpuregs_29_[4]), .B(_2104__bF_buf7), .Y(_2109_) );
OAI21X1 OAI21X1_2845 ( .A(_4955__bF_buf0), .B(_2104__bF_buf6), .C(_2109_), .Y(_447_) );
NAND2X1 NAND2X1_899 ( .A(cpuregs_29_[5]), .B(_2104__bF_buf5), .Y(_2110_) );
OAI21X1 OAI21X1_2846 ( .A(_4654__bF_buf4), .B(_2104__bF_buf4), .C(_2110_), .Y(_448_) );
NAND2X1 NAND2X1_900 ( .A(cpuregs_29_[6]), .B(_2104__bF_buf3), .Y(_2111_) );
OAI21X1 OAI21X1_2847 ( .A(_4664__bF_buf4), .B(_2104__bF_buf2), .C(_2111_), .Y(_449_) );
NAND2X1 NAND2X1_901 ( .A(cpuregs_29_[7]), .B(_2104__bF_buf1), .Y(_2112_) );
OAI21X1 OAI21X1_2848 ( .A(_4677__bF_buf4), .B(_2104__bF_buf0), .C(_2112_), .Y(_450_) );
NAND2X1 NAND2X1_902 ( .A(cpuregs_29_[8]), .B(_2104__bF_buf7), .Y(_2113_) );
OAI21X1 OAI21X1_2849 ( .A(_4685__bF_buf4), .B(_2104__bF_buf6), .C(_2113_), .Y(_451_) );
NAND2X1 NAND2X1_903 ( .A(cpuregs_29_[9]), .B(_2104__bF_buf5), .Y(_2114_) );
OAI21X1 OAI21X1_2850 ( .A(_4696__bF_buf4), .B(_2104__bF_buf4), .C(_2114_), .Y(_452_) );
NAND2X1 NAND2X1_904 ( .A(cpuregs_29_[10]), .B(_2104__bF_buf3), .Y(_2115_) );
OAI21X1 OAI21X1_2851 ( .A(_4703__bF_buf4), .B(_2104__bF_buf2), .C(_2115_), .Y(_453_) );
NAND2X1 NAND2X1_905 ( .A(cpuregs_29_[11]), .B(_2104__bF_buf1), .Y(_2116_) );
OAI21X1 OAI21X1_2852 ( .A(_4713__bF_buf4), .B(_2104__bF_buf0), .C(_2116_), .Y(_454_) );
NAND2X1 NAND2X1_906 ( .A(cpuregs_29_[12]), .B(_2104__bF_buf7), .Y(_2117_) );
OAI21X1 OAI21X1_2853 ( .A(_4722__bF_buf4), .B(_2104__bF_buf6), .C(_2117_), .Y(_455_) );
NAND2X1 NAND2X1_907 ( .A(cpuregs_29_[13]), .B(_2104__bF_buf5), .Y(_2118_) );
OAI21X1 OAI21X1_2854 ( .A(_4731__bF_buf4), .B(_2104__bF_buf4), .C(_2118_), .Y(_456_) );
NAND2X1 NAND2X1_908 ( .A(cpuregs_29_[14]), .B(_2104__bF_buf3), .Y(_2119_) );
OAI21X1 OAI21X1_2855 ( .A(_4740__bF_buf4), .B(_2104__bF_buf2), .C(_2119_), .Y(_457_) );
NAND2X1 NAND2X1_909 ( .A(cpuregs_29_[15]), .B(_2104__bF_buf1), .Y(_2120_) );
OAI21X1 OAI21X1_2856 ( .A(_4747__bF_buf4), .B(_2104__bF_buf0), .C(_2120_), .Y(_458_) );
NAND2X1 NAND2X1_910 ( .A(cpuregs_29_[16]), .B(_2104__bF_buf7), .Y(_2121_) );
OAI21X1 OAI21X1_2857 ( .A(_4755__bF_buf4), .B(_2104__bF_buf6), .C(_2121_), .Y(_459_) );
NAND2X1 NAND2X1_911 ( .A(cpuregs_29_[17]), .B(_2104__bF_buf5), .Y(_2122_) );
OAI21X1 OAI21X1_2858 ( .A(_4763__bF_buf4), .B(_2104__bF_buf4), .C(_2122_), .Y(_460_) );
NAND2X1 NAND2X1_912 ( .A(cpuregs_29_[18]), .B(_2104__bF_buf3), .Y(_2123_) );
OAI21X1 OAI21X1_2859 ( .A(_4783__bF_buf4), .B(_2104__bF_buf2), .C(_2123_), .Y(_461_) );
NAND2X1 NAND2X1_913 ( .A(cpuregs_29_[19]), .B(_2104__bF_buf1), .Y(_2124_) );
OAI21X1 OAI21X1_2860 ( .A(_4793__bF_buf4), .B(_2104__bF_buf0), .C(_2124_), .Y(_462_) );
NAND2X1 NAND2X1_914 ( .A(cpuregs_29_[20]), .B(_2104__bF_buf7), .Y(_2125_) );
OAI21X1 OAI21X1_2861 ( .A(_4806__bF_buf4), .B(_2104__bF_buf6), .C(_2125_), .Y(_463_) );
NAND2X1 NAND2X1_915 ( .A(cpuregs_29_[21]), .B(_2104__bF_buf5), .Y(_2126_) );
OAI21X1 OAI21X1_2862 ( .A(_4816__bF_buf4), .B(_2104__bF_buf4), .C(_2126_), .Y(_464_) );
NAND2X1 NAND2X1_916 ( .A(cpuregs_29_[22]), .B(_2104__bF_buf3), .Y(_2127_) );
OAI21X1 OAI21X1_2863 ( .A(_4824__bF_buf4), .B(_2104__bF_buf2), .C(_2127_), .Y(_465_) );
NAND2X1 NAND2X1_917 ( .A(cpuregs_29_[23]), .B(_2104__bF_buf1), .Y(_2128_) );
OAI21X1 OAI21X1_2864 ( .A(_4833__bF_buf4), .B(_2104__bF_buf0), .C(_2128_), .Y(_466_) );
NAND2X1 NAND2X1_918 ( .A(cpuregs_29_[24]), .B(_2104__bF_buf7), .Y(_2129_) );
OAI21X1 OAI21X1_2865 ( .A(_4845__bF_buf4), .B(_2104__bF_buf6), .C(_2129_), .Y(_467_) );
NAND2X1 NAND2X1_919 ( .A(cpuregs_29_[25]), .B(_2104__bF_buf5), .Y(_2130_) );
OAI21X1 OAI21X1_2866 ( .A(_4854__bF_buf4), .B(_2104__bF_buf4), .C(_2130_), .Y(_468_) );
NAND2X1 NAND2X1_920 ( .A(cpuregs_29_[26]), .B(_2104__bF_buf3), .Y(_2131_) );
OAI21X1 OAI21X1_2867 ( .A(_4863__bF_buf4), .B(_2104__bF_buf2), .C(_2131_), .Y(_469_) );
NAND2X1 NAND2X1_921 ( .A(cpuregs_29_[27]), .B(_2104__bF_buf1), .Y(_2132_) );
OAI21X1 OAI21X1_2868 ( .A(_4871__bF_buf4), .B(_2104__bF_buf0), .C(_2132_), .Y(_470_) );
NAND2X1 NAND2X1_922 ( .A(cpuregs_29_[28]), .B(_2104__bF_buf7), .Y(_2133_) );
OAI21X1 OAI21X1_2869 ( .A(_4884__bF_buf4), .B(_2104__bF_buf6), .C(_2133_), .Y(_471_) );
NAND2X1 NAND2X1_923 ( .A(cpuregs_29_[29]), .B(_2104__bF_buf5), .Y(_2134_) );
OAI21X1 OAI21X1_2870 ( .A(_4893__bF_buf4), .B(_2104__bF_buf4), .C(_2134_), .Y(_472_) );
NAND2X1 NAND2X1_924 ( .A(cpuregs_29_[30]), .B(_2104__bF_buf3), .Y(_2135_) );
OAI21X1 OAI21X1_2871 ( .A(_4901__bF_buf4), .B(_2104__bF_buf2), .C(_2135_), .Y(_473_) );
NAND2X1 NAND2X1_925 ( .A(cpuregs_29_[31]), .B(_2104__bF_buf1), .Y(_2136_) );
OAI21X1 OAI21X1_2872 ( .A(_4910__bF_buf4), .B(_2104__bF_buf0), .C(_2136_), .Y(_474_) );
NOR2X1 NOR2X1_1219 ( .A(_2035__bF_buf5), .B(_5706__bF_buf2), .Y(_2137_) );
INVX1 INVX1_1174 ( .A(_2137_), .Y(_2138_) );
OAI21X1 OAI21X1_2873 ( .A(_5706__bF_buf1), .B(_2035__bF_buf4), .C(cpuregs_28_[0]), .Y(_2139_) );
OAI21X1 OAI21X1_2874 ( .A(_2138__bF_buf4), .B(_4925__bF_buf4), .C(_2139_), .Y(_475_) );
OAI21X1 OAI21X1_2875 ( .A(_5706__bF_buf0), .B(_2035__bF_buf3), .C(cpuregs_28_[1]), .Y(_2140_) );
OAI21X1 OAI21X1_2876 ( .A(_2138__bF_buf3), .B(_4933__bF_buf4), .C(_2140_), .Y(_476_) );
OAI21X1 OAI21X1_2877 ( .A(_5706__bF_buf11), .B(_2035__bF_buf2), .C(cpuregs_28_[2]), .Y(_2141_) );
OAI21X1 OAI21X1_2878 ( .A(_2138__bF_buf2), .B(_4940__bF_buf4), .C(_2141_), .Y(_477_) );
OAI21X1 OAI21X1_2879 ( .A(_5706__bF_buf10), .B(_2035__bF_buf1), .C(cpuregs_28_[3]), .Y(_2142_) );
OAI21X1 OAI21X1_2880 ( .A(_2138__bF_buf1), .B(_4948__bF_buf4), .C(_2142_), .Y(_478_) );
OAI21X1 OAI21X1_2881 ( .A(_5706__bF_buf9), .B(_2035__bF_buf0), .C(cpuregs_28_[4]), .Y(_2143_) );
OAI21X1 OAI21X1_2882 ( .A(_2138__bF_buf0), .B(_4955__bF_buf4), .C(_2143_), .Y(_479_) );
OAI21X1 OAI21X1_2883 ( .A(_5706__bF_buf8), .B(_2035__bF_buf8), .C(cpuregs_28_[5]), .Y(_2144_) );
OAI21X1 OAI21X1_2884 ( .A(_2138__bF_buf4), .B(_4654__bF_buf3), .C(_2144_), .Y(_480_) );
OAI21X1 OAI21X1_2885 ( .A(_5706__bF_buf7), .B(_2035__bF_buf7), .C(cpuregs_28_[6]), .Y(_2145_) );
OAI21X1 OAI21X1_2886 ( .A(_2138__bF_buf3), .B(_4664__bF_buf3), .C(_2145_), .Y(_481_) );
OAI21X1 OAI21X1_2887 ( .A(_5706__bF_buf6), .B(_2035__bF_buf6), .C(cpuregs_28_[7]), .Y(_2146_) );
OAI21X1 OAI21X1_2888 ( .A(_2138__bF_buf2), .B(_4677__bF_buf3), .C(_2146_), .Y(_482_) );
OAI21X1 OAI21X1_2889 ( .A(_5706__bF_buf5), .B(_2035__bF_buf5), .C(cpuregs_28_[8]), .Y(_2147_) );
OAI21X1 OAI21X1_2890 ( .A(_4685__bF_buf3), .B(_2138__bF_buf1), .C(_2147_), .Y(_483_) );
OAI21X1 OAI21X1_2891 ( .A(_5706__bF_buf4), .B(_2035__bF_buf4), .C(cpuregs_28_[9]), .Y(_2148_) );
OAI21X1 OAI21X1_2892 ( .A(_4696__bF_buf3), .B(_2138__bF_buf0), .C(_2148_), .Y(_484_) );
OAI21X1 OAI21X1_2893 ( .A(_5706__bF_buf3), .B(_2035__bF_buf3), .C(cpuregs_28_[10]), .Y(_2149_) );
OAI21X1 OAI21X1_2894 ( .A(_4703__bF_buf3), .B(_2138__bF_buf4), .C(_2149_), .Y(_485_) );
OAI21X1 OAI21X1_2895 ( .A(_5706__bF_buf2), .B(_2035__bF_buf2), .C(cpuregs_28_[11]), .Y(_2150_) );
OAI21X1 OAI21X1_2896 ( .A(_4713__bF_buf3), .B(_2138__bF_buf3), .C(_2150_), .Y(_486_) );
OAI21X1 OAI21X1_2897 ( .A(_5706__bF_buf1), .B(_2035__bF_buf1), .C(cpuregs_28_[12]), .Y(_2151_) );
OAI21X1 OAI21X1_2898 ( .A(_4722__bF_buf3), .B(_2138__bF_buf2), .C(_2151_), .Y(_487_) );
OAI21X1 OAI21X1_2899 ( .A(_5706__bF_buf0), .B(_2035__bF_buf0), .C(cpuregs_28_[13]), .Y(_2152_) );
OAI21X1 OAI21X1_2900 ( .A(_4731__bF_buf3), .B(_2138__bF_buf1), .C(_2152_), .Y(_488_) );
OAI21X1 OAI21X1_2901 ( .A(_5706__bF_buf11), .B(_2035__bF_buf8), .C(cpuregs_28_[14]), .Y(_2153_) );
OAI21X1 OAI21X1_2902 ( .A(_4740__bF_buf3), .B(_2138__bF_buf0), .C(_2153_), .Y(_489_) );
OAI21X1 OAI21X1_2903 ( .A(_5706__bF_buf10), .B(_2035__bF_buf7), .C(cpuregs_28_[15]), .Y(_2154_) );
OAI21X1 OAI21X1_2904 ( .A(_4747__bF_buf3), .B(_2138__bF_buf4), .C(_2154_), .Y(_490_) );
OAI21X1 OAI21X1_2905 ( .A(_5706__bF_buf9), .B(_2035__bF_buf6), .C(cpuregs_28_[16]), .Y(_2155_) );
OAI21X1 OAI21X1_2906 ( .A(_4755__bF_buf3), .B(_2138__bF_buf3), .C(_2155_), .Y(_491_) );
OAI21X1 OAI21X1_2907 ( .A(_5706__bF_buf8), .B(_2035__bF_buf5), .C(cpuregs_28_[17]), .Y(_2156_) );
OAI21X1 OAI21X1_2908 ( .A(_4763__bF_buf3), .B(_2138__bF_buf2), .C(_2156_), .Y(_492_) );
OAI21X1 OAI21X1_2909 ( .A(_5706__bF_buf7), .B(_2035__bF_buf4), .C(cpuregs_28_[18]), .Y(_2157_) );
OAI21X1 OAI21X1_2910 ( .A(_4783__bF_buf3), .B(_2138__bF_buf1), .C(_2157_), .Y(_493_) );
OAI21X1 OAI21X1_2911 ( .A(_5706__bF_buf6), .B(_2035__bF_buf3), .C(cpuregs_28_[19]), .Y(_2158_) );
OAI21X1 OAI21X1_2912 ( .A(_4793__bF_buf3), .B(_2138__bF_buf0), .C(_2158_), .Y(_494_) );
OAI21X1 OAI21X1_2913 ( .A(_5706__bF_buf5), .B(_2035__bF_buf2), .C(cpuregs_28_[20]), .Y(_2159_) );
OAI21X1 OAI21X1_2914 ( .A(_4806__bF_buf3), .B(_2138__bF_buf4), .C(_2159_), .Y(_495_) );
OAI21X1 OAI21X1_2915 ( .A(_5706__bF_buf4), .B(_2035__bF_buf1), .C(cpuregs_28_[21]), .Y(_2160_) );
OAI21X1 OAI21X1_2916 ( .A(_4816__bF_buf3), .B(_2138__bF_buf3), .C(_2160_), .Y(_496_) );
OAI21X1 OAI21X1_2917 ( .A(_5706__bF_buf3), .B(_2035__bF_buf0), .C(cpuregs_28_[22]), .Y(_2161_) );
OAI21X1 OAI21X1_2918 ( .A(_4824__bF_buf3), .B(_2138__bF_buf2), .C(_2161_), .Y(_497_) );
OAI21X1 OAI21X1_2919 ( .A(_5706__bF_buf2), .B(_2035__bF_buf8), .C(cpuregs_28_[23]), .Y(_2162_) );
OAI21X1 OAI21X1_2920 ( .A(_4833__bF_buf3), .B(_2138__bF_buf1), .C(_2162_), .Y(_498_) );
OAI21X1 OAI21X1_2921 ( .A(_5706__bF_buf1), .B(_2035__bF_buf7), .C(cpuregs_28_[24]), .Y(_2163_) );
OAI21X1 OAI21X1_2922 ( .A(_4845__bF_buf3), .B(_2138__bF_buf0), .C(_2163_), .Y(_499_) );
OAI21X1 OAI21X1_2923 ( .A(_5706__bF_buf0), .B(_2035__bF_buf6), .C(cpuregs_28_[25]), .Y(_2164_) );
OAI21X1 OAI21X1_2924 ( .A(_4854__bF_buf3), .B(_2138__bF_buf4), .C(_2164_), .Y(_500_) );
OAI21X1 OAI21X1_2925 ( .A(_5706__bF_buf11), .B(_2035__bF_buf5), .C(cpuregs_28_[26]), .Y(_2165_) );
OAI21X1 OAI21X1_2926 ( .A(_4863__bF_buf3), .B(_2138__bF_buf3), .C(_2165_), .Y(_501_) );
OAI21X1 OAI21X1_2927 ( .A(_5706__bF_buf10), .B(_2035__bF_buf4), .C(cpuregs_28_[27]), .Y(_2166_) );
OAI21X1 OAI21X1_2928 ( .A(_4871__bF_buf3), .B(_2138__bF_buf2), .C(_2166_), .Y(_502_) );
OAI21X1 OAI21X1_2929 ( .A(_5706__bF_buf9), .B(_2035__bF_buf3), .C(cpuregs_28_[28]), .Y(_2167_) );
OAI21X1 OAI21X1_2930 ( .A(_4884__bF_buf3), .B(_2138__bF_buf1), .C(_2167_), .Y(_503_) );
OAI21X1 OAI21X1_2931 ( .A(_5706__bF_buf8), .B(_2035__bF_buf2), .C(cpuregs_28_[29]), .Y(_2168_) );
OAI21X1 OAI21X1_2932 ( .A(_4893__bF_buf3), .B(_2138__bF_buf0), .C(_2168_), .Y(_504_) );
OAI21X1 OAI21X1_2933 ( .A(_5706__bF_buf7), .B(_2035__bF_buf1), .C(cpuregs_28_[30]), .Y(_2169_) );
OAI21X1 OAI21X1_2934 ( .A(_4901__bF_buf3), .B(_2138__bF_buf4), .C(_2169_), .Y(_505_) );
OAI21X1 OAI21X1_2935 ( .A(_5706__bF_buf6), .B(_2035__bF_buf0), .C(cpuregs_28_[31]), .Y(_2170_) );
OAI21X1 OAI21X1_2936 ( .A(_4910__bF_buf3), .B(_2138__bF_buf3), .C(_2170_), .Y(_506_) );
NAND2X1 NAND2X1_926 ( .A(_4911_), .B(_2034_), .Y(_2171_) );
NOR2X1 NOR2X1_1220 ( .A(_2171__bF_buf8), .B(_4917__bF_buf10), .Y(_2172_) );
INVX1 INVX1_1175 ( .A(_2172_), .Y(_2173_) );
OAI21X1 OAI21X1_2937 ( .A(_4917__bF_buf9), .B(_2171__bF_buf7), .C(cpuregs_27_[0]), .Y(_2174_) );
OAI21X1 OAI21X1_2938 ( .A(_2173__bF_buf4), .B(_4925__bF_buf3), .C(_2174_), .Y(_507_) );
OAI21X1 OAI21X1_2939 ( .A(_4917__bF_buf8), .B(_2171__bF_buf6), .C(cpuregs_27_[1]), .Y(_2175_) );
OAI21X1 OAI21X1_2940 ( .A(_2173__bF_buf3), .B(_4933__bF_buf3), .C(_2175_), .Y(_508_) );
OAI21X1 OAI21X1_2941 ( .A(_4917__bF_buf7), .B(_2171__bF_buf5), .C(cpuregs_27_[2]), .Y(_2176_) );
OAI21X1 OAI21X1_2942 ( .A(_2173__bF_buf2), .B(_4940__bF_buf3), .C(_2176_), .Y(_509_) );
OAI21X1 OAI21X1_2943 ( .A(_4917__bF_buf6), .B(_2171__bF_buf4), .C(cpuregs_27_[3]), .Y(_2177_) );
OAI21X1 OAI21X1_2944 ( .A(_2173__bF_buf1), .B(_4948__bF_buf3), .C(_2177_), .Y(_510_) );
OAI21X1 OAI21X1_2945 ( .A(_4917__bF_buf5), .B(_2171__bF_buf3), .C(cpuregs_27_[4]), .Y(_2178_) );
OAI21X1 OAI21X1_2946 ( .A(_2173__bF_buf0), .B(_4955__bF_buf3), .C(_2178_), .Y(_511_) );
OAI21X1 OAI21X1_2947 ( .A(_4917__bF_buf4), .B(_2171__bF_buf2), .C(cpuregs_27_[5]), .Y(_2179_) );
OAI21X1 OAI21X1_2948 ( .A(_2173__bF_buf4), .B(_4654__bF_buf2), .C(_2179_), .Y(_512_) );
OAI21X1 OAI21X1_2949 ( .A(_4917__bF_buf3), .B(_2171__bF_buf1), .C(cpuregs_27_[6]), .Y(_2180_) );
OAI21X1 OAI21X1_2950 ( .A(_4664__bF_buf2), .B(_2173__bF_buf3), .C(_2180_), .Y(_513_) );
OAI21X1 OAI21X1_2951 ( .A(_4917__bF_buf2), .B(_2171__bF_buf0), .C(cpuregs_27_[7]), .Y(_2181_) );
OAI21X1 OAI21X1_2952 ( .A(_4677__bF_buf2), .B(_2173__bF_buf2), .C(_2181_), .Y(_514_) );
OAI21X1 OAI21X1_2953 ( .A(_4917__bF_buf1), .B(_2171__bF_buf8), .C(cpuregs_27_[8]), .Y(_2182_) );
OAI21X1 OAI21X1_2954 ( .A(_4685__bF_buf2), .B(_2173__bF_buf1), .C(_2182_), .Y(_515_) );
OAI21X1 OAI21X1_2955 ( .A(_4917__bF_buf0), .B(_2171__bF_buf7), .C(cpuregs_27_[9]), .Y(_2183_) );
OAI21X1 OAI21X1_2956 ( .A(_4696__bF_buf2), .B(_2173__bF_buf0), .C(_2183_), .Y(_516_) );
OAI21X1 OAI21X1_2957 ( .A(_4917__bF_buf10), .B(_2171__bF_buf6), .C(cpuregs_27_[10]), .Y(_2184_) );
OAI21X1 OAI21X1_2958 ( .A(_4703__bF_buf2), .B(_2173__bF_buf4), .C(_2184_), .Y(_517_) );
OAI21X1 OAI21X1_2959 ( .A(_4917__bF_buf9), .B(_2171__bF_buf5), .C(cpuregs_27_[11]), .Y(_2185_) );
OAI21X1 OAI21X1_2960 ( .A(_4713__bF_buf2), .B(_2173__bF_buf3), .C(_2185_), .Y(_518_) );
OAI21X1 OAI21X1_2961 ( .A(_4917__bF_buf8), .B(_2171__bF_buf4), .C(cpuregs_27_[12]), .Y(_2186_) );
OAI21X1 OAI21X1_2962 ( .A(_4722__bF_buf2), .B(_2173__bF_buf2), .C(_2186_), .Y(_519_) );
OAI21X1 OAI21X1_2963 ( .A(_4917__bF_buf7), .B(_2171__bF_buf3), .C(cpuregs_27_[13]), .Y(_2187_) );
OAI21X1 OAI21X1_2964 ( .A(_4731__bF_buf2), .B(_2173__bF_buf1), .C(_2187_), .Y(_520_) );
OAI21X1 OAI21X1_2965 ( .A(_4917__bF_buf6), .B(_2171__bF_buf2), .C(cpuregs_27_[14]), .Y(_2188_) );
OAI21X1 OAI21X1_2966 ( .A(_4740__bF_buf2), .B(_2173__bF_buf0), .C(_2188_), .Y(_521_) );
OAI21X1 OAI21X1_2967 ( .A(_4917__bF_buf5), .B(_2171__bF_buf1), .C(cpuregs_27_[15]), .Y(_2189_) );
OAI21X1 OAI21X1_2968 ( .A(_4747__bF_buf2), .B(_2173__bF_buf4), .C(_2189_), .Y(_522_) );
OAI21X1 OAI21X1_2969 ( .A(_4917__bF_buf4), .B(_2171__bF_buf0), .C(cpuregs_27_[16]), .Y(_2190_) );
OAI21X1 OAI21X1_2970 ( .A(_4755__bF_buf2), .B(_2173__bF_buf3), .C(_2190_), .Y(_523_) );
OAI21X1 OAI21X1_2971 ( .A(_4917__bF_buf3), .B(_2171__bF_buf8), .C(cpuregs_27_[17]), .Y(_2191_) );
OAI21X1 OAI21X1_2972 ( .A(_4763__bF_buf2), .B(_2173__bF_buf2), .C(_2191_), .Y(_524_) );
OAI21X1 OAI21X1_2973 ( .A(_4917__bF_buf2), .B(_2171__bF_buf7), .C(cpuregs_27_[18]), .Y(_2192_) );
OAI21X1 OAI21X1_2974 ( .A(_4783__bF_buf2), .B(_2173__bF_buf1), .C(_2192_), .Y(_525_) );
OAI21X1 OAI21X1_2975 ( .A(_4917__bF_buf1), .B(_2171__bF_buf6), .C(cpuregs_27_[19]), .Y(_2193_) );
OAI21X1 OAI21X1_2976 ( .A(_4793__bF_buf2), .B(_2173__bF_buf0), .C(_2193_), .Y(_526_) );
OAI21X1 OAI21X1_2977 ( .A(_4917__bF_buf0), .B(_2171__bF_buf5), .C(cpuregs_27_[20]), .Y(_2194_) );
OAI21X1 OAI21X1_2978 ( .A(_4806__bF_buf2), .B(_2173__bF_buf4), .C(_2194_), .Y(_527_) );
OAI21X1 OAI21X1_2979 ( .A(_4917__bF_buf10), .B(_2171__bF_buf4), .C(cpuregs_27_[21]), .Y(_2195_) );
OAI21X1 OAI21X1_2980 ( .A(_4816__bF_buf2), .B(_2173__bF_buf3), .C(_2195_), .Y(_528_) );
OAI21X1 OAI21X1_2981 ( .A(_4917__bF_buf9), .B(_2171__bF_buf3), .C(cpuregs_27_[22]), .Y(_2196_) );
OAI21X1 OAI21X1_2982 ( .A(_4824__bF_buf2), .B(_2173__bF_buf2), .C(_2196_), .Y(_529_) );
OAI21X1 OAI21X1_2983 ( .A(_4917__bF_buf8), .B(_2171__bF_buf2), .C(cpuregs_27_[23]), .Y(_2197_) );
OAI21X1 OAI21X1_2984 ( .A(_4833__bF_buf2), .B(_2173__bF_buf1), .C(_2197_), .Y(_530_) );
OAI21X1 OAI21X1_2985 ( .A(_4917__bF_buf7), .B(_2171__bF_buf1), .C(cpuregs_27_[24]), .Y(_2198_) );
OAI21X1 OAI21X1_2986 ( .A(_4845__bF_buf2), .B(_2173__bF_buf0), .C(_2198_), .Y(_531_) );
OAI21X1 OAI21X1_2987 ( .A(_4917__bF_buf6), .B(_2171__bF_buf0), .C(cpuregs_27_[25]), .Y(_2199_) );
OAI21X1 OAI21X1_2988 ( .A(_4854__bF_buf2), .B(_2173__bF_buf4), .C(_2199_), .Y(_532_) );
OAI21X1 OAI21X1_2989 ( .A(_4917__bF_buf5), .B(_2171__bF_buf8), .C(cpuregs_27_[26]), .Y(_2200_) );
OAI21X1 OAI21X1_2990 ( .A(_4863__bF_buf2), .B(_2173__bF_buf3), .C(_2200_), .Y(_533_) );
OAI21X1 OAI21X1_2991 ( .A(_4917__bF_buf4), .B(_2171__bF_buf7), .C(cpuregs_27_[27]), .Y(_2201_) );
OAI21X1 OAI21X1_2992 ( .A(_4871__bF_buf2), .B(_2173__bF_buf2), .C(_2201_), .Y(_534_) );
OAI21X1 OAI21X1_2993 ( .A(_4917__bF_buf3), .B(_2171__bF_buf6), .C(cpuregs_27_[28]), .Y(_2202_) );
OAI21X1 OAI21X1_2994 ( .A(_4884__bF_buf2), .B(_2173__bF_buf1), .C(_2202_), .Y(_535_) );
OAI21X1 OAI21X1_2995 ( .A(_4917__bF_buf2), .B(_2171__bF_buf5), .C(cpuregs_27_[29]), .Y(_2203_) );
OAI21X1 OAI21X1_2996 ( .A(_4893__bF_buf2), .B(_2173__bF_buf0), .C(_2203_), .Y(_536_) );
OAI21X1 OAI21X1_2997 ( .A(_4917__bF_buf1), .B(_2171__bF_buf4), .C(cpuregs_27_[30]), .Y(_2204_) );
OAI21X1 OAI21X1_2998 ( .A(_4901__bF_buf2), .B(_2173__bF_buf4), .C(_2204_), .Y(_537_) );
OAI21X1 OAI21X1_2999 ( .A(_4917__bF_buf0), .B(_2171__bF_buf3), .C(cpuregs_27_[31]), .Y(_2205_) );
OAI21X1 OAI21X1_3000 ( .A(_4910__bF_buf2), .B(_2173__bF_buf3), .C(_2205_), .Y(_538_) );
NOR2X1 NOR2X1_1221 ( .A(_2171__bF_buf2), .B(_5281__bF_buf8), .Y(_2206_) );
INVX1 INVX1_1176 ( .A(_2206_), .Y(_2207_) );
OAI21X1 OAI21X1_3001 ( .A(_5281__bF_buf7), .B(_2171__bF_buf1), .C(cpuregs_26_[0]), .Y(_2208_) );
OAI21X1 OAI21X1_3002 ( .A(_2207__bF_buf4), .B(_4925__bF_buf2), .C(_2208_), .Y(_539_) );
OAI21X1 OAI21X1_3003 ( .A(_5281__bF_buf6), .B(_2171__bF_buf0), .C(cpuregs_26_[1]), .Y(_2209_) );
OAI21X1 OAI21X1_3004 ( .A(_2207__bF_buf3), .B(_4933__bF_buf2), .C(_2209_), .Y(_540_) );
OAI21X1 OAI21X1_3005 ( .A(_5281__bF_buf5), .B(_2171__bF_buf8), .C(cpuregs_26_[2]), .Y(_2210_) );
OAI21X1 OAI21X1_3006 ( .A(_2207__bF_buf2), .B(_4940__bF_buf2), .C(_2210_), .Y(_541_) );
OAI21X1 OAI21X1_3007 ( .A(_5281__bF_buf4), .B(_2171__bF_buf7), .C(cpuregs_26_[3]), .Y(_2211_) );
OAI21X1 OAI21X1_3008 ( .A(_2207__bF_buf1), .B(_4948__bF_buf2), .C(_2211_), .Y(_542_) );
OAI21X1 OAI21X1_3009 ( .A(_5281__bF_buf3), .B(_2171__bF_buf6), .C(cpuregs_26_[4]), .Y(_2212_) );
OAI21X1 OAI21X1_3010 ( .A(_2207__bF_buf0), .B(_4955__bF_buf2), .C(_2212_), .Y(_543_) );
OAI21X1 OAI21X1_3011 ( .A(_5281__bF_buf2), .B(_2171__bF_buf5), .C(cpuregs_26_[5]), .Y(_2213_) );
OAI21X1 OAI21X1_3012 ( .A(_2207__bF_buf4), .B(_4654__bF_buf1), .C(_2213_), .Y(_544_) );
OAI21X1 OAI21X1_3013 ( .A(_5281__bF_buf1), .B(_2171__bF_buf4), .C(cpuregs_26_[6]), .Y(_2214_) );
OAI21X1 OAI21X1_3014 ( .A(_4664__bF_buf1), .B(_2207__bF_buf3), .C(_2214_), .Y(_545_) );
OAI21X1 OAI21X1_3015 ( .A(_5281__bF_buf0), .B(_2171__bF_buf3), .C(cpuregs_26_[7]), .Y(_2215_) );
OAI21X1 OAI21X1_3016 ( .A(_4677__bF_buf1), .B(_2207__bF_buf2), .C(_2215_), .Y(_546_) );
OAI21X1 OAI21X1_3017 ( .A(_5281__bF_buf10), .B(_2171__bF_buf2), .C(cpuregs_26_[8]), .Y(_2216_) );
OAI21X1 OAI21X1_3018 ( .A(_4685__bF_buf1), .B(_2207__bF_buf1), .C(_2216_), .Y(_547_) );
OAI21X1 OAI21X1_3019 ( .A(_5281__bF_buf9), .B(_2171__bF_buf1), .C(cpuregs_26_[9]), .Y(_2217_) );
OAI21X1 OAI21X1_3020 ( .A(_4696__bF_buf1), .B(_2207__bF_buf0), .C(_2217_), .Y(_548_) );
OAI21X1 OAI21X1_3021 ( .A(_5281__bF_buf8), .B(_2171__bF_buf0), .C(cpuregs_26_[10]), .Y(_2218_) );
OAI21X1 OAI21X1_3022 ( .A(_4703__bF_buf1), .B(_2207__bF_buf4), .C(_2218_), .Y(_549_) );
OAI21X1 OAI21X1_3023 ( .A(_5281__bF_buf7), .B(_2171__bF_buf8), .C(cpuregs_26_[11]), .Y(_2219_) );
OAI21X1 OAI21X1_3024 ( .A(_4713__bF_buf1), .B(_2207__bF_buf3), .C(_2219_), .Y(_550_) );
OAI21X1 OAI21X1_3025 ( .A(_5281__bF_buf6), .B(_2171__bF_buf7), .C(cpuregs_26_[12]), .Y(_2220_) );
OAI21X1 OAI21X1_3026 ( .A(_4722__bF_buf1), .B(_2207__bF_buf2), .C(_2220_), .Y(_551_) );
OAI21X1 OAI21X1_3027 ( .A(_5281__bF_buf5), .B(_2171__bF_buf6), .C(cpuregs_26_[13]), .Y(_2221_) );
OAI21X1 OAI21X1_3028 ( .A(_4731__bF_buf1), .B(_2207__bF_buf1), .C(_2221_), .Y(_552_) );
OAI21X1 OAI21X1_3029 ( .A(_5281__bF_buf4), .B(_2171__bF_buf5), .C(cpuregs_26_[14]), .Y(_2222_) );
OAI21X1 OAI21X1_3030 ( .A(_4740__bF_buf1), .B(_2207__bF_buf0), .C(_2222_), .Y(_553_) );
OAI21X1 OAI21X1_3031 ( .A(_5281__bF_buf3), .B(_2171__bF_buf4), .C(cpuregs_26_[15]), .Y(_2223_) );
OAI21X1 OAI21X1_3032 ( .A(_4747__bF_buf1), .B(_2207__bF_buf4), .C(_2223_), .Y(_554_) );
OAI21X1 OAI21X1_3033 ( .A(_5281__bF_buf2), .B(_2171__bF_buf3), .C(cpuregs_26_[16]), .Y(_2224_) );
OAI21X1 OAI21X1_3034 ( .A(_4755__bF_buf1), .B(_2207__bF_buf3), .C(_2224_), .Y(_555_) );
OAI21X1 OAI21X1_3035 ( .A(_5281__bF_buf1), .B(_2171__bF_buf2), .C(cpuregs_26_[17]), .Y(_2225_) );
OAI21X1 OAI21X1_3036 ( .A(_4763__bF_buf1), .B(_2207__bF_buf2), .C(_2225_), .Y(_556_) );
OAI21X1 OAI21X1_3037 ( .A(_5281__bF_buf0), .B(_2171__bF_buf1), .C(cpuregs_26_[18]), .Y(_2226_) );
OAI21X1 OAI21X1_3038 ( .A(_4783__bF_buf1), .B(_2207__bF_buf1), .C(_2226_), .Y(_557_) );
OAI21X1 OAI21X1_3039 ( .A(_5281__bF_buf10), .B(_2171__bF_buf0), .C(cpuregs_26_[19]), .Y(_2227_) );
OAI21X1 OAI21X1_3040 ( .A(_4793__bF_buf1), .B(_2207__bF_buf0), .C(_2227_), .Y(_558_) );
OAI21X1 OAI21X1_3041 ( .A(_5281__bF_buf9), .B(_2171__bF_buf8), .C(cpuregs_26_[20]), .Y(_2228_) );
OAI21X1 OAI21X1_3042 ( .A(_4806__bF_buf1), .B(_2207__bF_buf4), .C(_2228_), .Y(_559_) );
OAI21X1 OAI21X1_3043 ( .A(_5281__bF_buf8), .B(_2171__bF_buf7), .C(cpuregs_26_[21]), .Y(_2229_) );
OAI21X1 OAI21X1_3044 ( .A(_4816__bF_buf1), .B(_2207__bF_buf3), .C(_2229_), .Y(_560_) );
OAI21X1 OAI21X1_3045 ( .A(_5281__bF_buf7), .B(_2171__bF_buf6), .C(cpuregs_26_[22]), .Y(_2230_) );
OAI21X1 OAI21X1_3046 ( .A(_4824__bF_buf1), .B(_2207__bF_buf2), .C(_2230_), .Y(_561_) );
OAI21X1 OAI21X1_3047 ( .A(_5281__bF_buf6), .B(_2171__bF_buf5), .C(cpuregs_26_[23]), .Y(_2231_) );
OAI21X1 OAI21X1_3048 ( .A(_4833__bF_buf1), .B(_2207__bF_buf1), .C(_2231_), .Y(_562_) );
OAI21X1 OAI21X1_3049 ( .A(_5281__bF_buf5), .B(_2171__bF_buf4), .C(cpuregs_26_[24]), .Y(_2232_) );
OAI21X1 OAI21X1_3050 ( .A(_4845__bF_buf1), .B(_2207__bF_buf0), .C(_2232_), .Y(_563_) );
OAI21X1 OAI21X1_3051 ( .A(_5281__bF_buf4), .B(_2171__bF_buf3), .C(cpuregs_26_[25]), .Y(_2233_) );
OAI21X1 OAI21X1_3052 ( .A(_4854__bF_buf1), .B(_2207__bF_buf4), .C(_2233_), .Y(_564_) );
OAI21X1 OAI21X1_3053 ( .A(_5281__bF_buf3), .B(_2171__bF_buf2), .C(cpuregs_26_[26]), .Y(_2234_) );
OAI21X1 OAI21X1_3054 ( .A(_4863__bF_buf1), .B(_2207__bF_buf3), .C(_2234_), .Y(_565_) );
OAI21X1 OAI21X1_3055 ( .A(_5281__bF_buf2), .B(_2171__bF_buf1), .C(cpuregs_26_[27]), .Y(_2235_) );
OAI21X1 OAI21X1_3056 ( .A(_4871__bF_buf1), .B(_2207__bF_buf2), .C(_2235_), .Y(_566_) );
OAI21X1 OAI21X1_3057 ( .A(_5281__bF_buf1), .B(_2171__bF_buf0), .C(cpuregs_26_[28]), .Y(_2236_) );
OAI21X1 OAI21X1_3058 ( .A(_4884__bF_buf1), .B(_2207__bF_buf1), .C(_2236_), .Y(_567_) );
OAI21X1 OAI21X1_3059 ( .A(_5281__bF_buf0), .B(_2171__bF_buf8), .C(cpuregs_26_[29]), .Y(_2237_) );
OAI21X1 OAI21X1_3060 ( .A(_4893__bF_buf1), .B(_2207__bF_buf0), .C(_2237_), .Y(_568_) );
OAI21X1 OAI21X1_3061 ( .A(_5281__bF_buf10), .B(_2171__bF_buf7), .C(cpuregs_26_[30]), .Y(_2238_) );
OAI21X1 OAI21X1_3062 ( .A(_4901__bF_buf1), .B(_2207__bF_buf4), .C(_2238_), .Y(_569_) );
OAI21X1 OAI21X1_3063 ( .A(_5281__bF_buf9), .B(_2171__bF_buf6), .C(cpuregs_26_[31]), .Y(_2239_) );
OAI21X1 OAI21X1_3064 ( .A(_4910__bF_buf1), .B(_2207__bF_buf3), .C(_2239_), .Y(_570_) );
NAND3X1 NAND3X1_93 ( .A(_4911_), .B(_2034_), .C(_5313_), .Y(_2240_) );
NAND2X1 NAND2X1_927 ( .A(cpuregs_25_[0]), .B(_2240__bF_buf7), .Y(_2241_) );
OAI21X1 OAI21X1_3065 ( .A(_4925__bF_buf1), .B(_2240__bF_buf6), .C(_2241_), .Y(_571_) );
NAND2X1 NAND2X1_928 ( .A(cpuregs_25_[1]), .B(_2240__bF_buf5), .Y(_2242_) );
OAI21X1 OAI21X1_3066 ( .A(_4933__bF_buf1), .B(_2240__bF_buf4), .C(_2242_), .Y(_572_) );
NAND2X1 NAND2X1_929 ( .A(cpuregs_25_[2]), .B(_2240__bF_buf3), .Y(_2243_) );
OAI21X1 OAI21X1_3067 ( .A(_4940__bF_buf1), .B(_2240__bF_buf2), .C(_2243_), .Y(_573_) );
NAND2X1 NAND2X1_930 ( .A(cpuregs_25_[3]), .B(_2240__bF_buf1), .Y(_2244_) );
OAI21X1 OAI21X1_3068 ( .A(_4948__bF_buf1), .B(_2240__bF_buf0), .C(_2244_), .Y(_574_) );
NAND2X1 NAND2X1_931 ( .A(cpuregs_25_[4]), .B(_2240__bF_buf7), .Y(_2245_) );
OAI21X1 OAI21X1_3069 ( .A(_4955__bF_buf1), .B(_2240__bF_buf6), .C(_2245_), .Y(_575_) );
NAND2X1 NAND2X1_932 ( .A(cpuregs_25_[5]), .B(_2240__bF_buf5), .Y(_2246_) );
OAI21X1 OAI21X1_3070 ( .A(_4654__bF_buf0), .B(_2240__bF_buf4), .C(_2246_), .Y(_576_) );
NAND2X1 NAND2X1_933 ( .A(cpuregs_25_[6]), .B(_2240__bF_buf3), .Y(_2247_) );
OAI21X1 OAI21X1_3071 ( .A(_4664__bF_buf0), .B(_2240__bF_buf2), .C(_2247_), .Y(_577_) );
NAND2X1 NAND2X1_934 ( .A(cpuregs_25_[7]), .B(_2240__bF_buf1), .Y(_2248_) );
OAI21X1 OAI21X1_3072 ( .A(_4677__bF_buf0), .B(_2240__bF_buf0), .C(_2248_), .Y(_578_) );
NAND2X1 NAND2X1_935 ( .A(cpuregs_25_[8]), .B(_2240__bF_buf7), .Y(_2249_) );
OAI21X1 OAI21X1_3073 ( .A(_4685__bF_buf0), .B(_2240__bF_buf6), .C(_2249_), .Y(_579_) );
NAND2X1 NAND2X1_936 ( .A(cpuregs_25_[9]), .B(_2240__bF_buf5), .Y(_2250_) );
OAI21X1 OAI21X1_3074 ( .A(_4696__bF_buf0), .B(_2240__bF_buf4), .C(_2250_), .Y(_580_) );
NAND2X1 NAND2X1_937 ( .A(cpuregs_25_[10]), .B(_2240__bF_buf3), .Y(_2251_) );
OAI21X1 OAI21X1_3075 ( .A(_4703__bF_buf0), .B(_2240__bF_buf2), .C(_2251_), .Y(_581_) );
NAND2X1 NAND2X1_938 ( .A(cpuregs_25_[11]), .B(_2240__bF_buf1), .Y(_2252_) );
OAI21X1 OAI21X1_3076 ( .A(_4713__bF_buf0), .B(_2240__bF_buf0), .C(_2252_), .Y(_582_) );
NAND2X1 NAND2X1_939 ( .A(cpuregs_25_[12]), .B(_2240__bF_buf7), .Y(_2253_) );
OAI21X1 OAI21X1_3077 ( .A(_4722__bF_buf0), .B(_2240__bF_buf6), .C(_2253_), .Y(_583_) );
NAND2X1 NAND2X1_940 ( .A(cpuregs_25_[13]), .B(_2240__bF_buf5), .Y(_2254_) );
OAI21X1 OAI21X1_3078 ( .A(_4731__bF_buf0), .B(_2240__bF_buf4), .C(_2254_), .Y(_584_) );
NAND2X1 NAND2X1_941 ( .A(cpuregs_25_[14]), .B(_2240__bF_buf3), .Y(_2255_) );
OAI21X1 OAI21X1_3079 ( .A(_4740__bF_buf0), .B(_2240__bF_buf2), .C(_2255_), .Y(_585_) );
NAND2X1 NAND2X1_942 ( .A(cpuregs_25_[15]), .B(_2240__bF_buf1), .Y(_2256_) );
OAI21X1 OAI21X1_3080 ( .A(_4747__bF_buf0), .B(_2240__bF_buf0), .C(_2256_), .Y(_586_) );
NAND2X1 NAND2X1_943 ( .A(cpuregs_25_[16]), .B(_2240__bF_buf7), .Y(_2257_) );
OAI21X1 OAI21X1_3081 ( .A(_4755__bF_buf0), .B(_2240__bF_buf6), .C(_2257_), .Y(_587_) );
NAND2X1 NAND2X1_944 ( .A(cpuregs_25_[17]), .B(_2240__bF_buf5), .Y(_2258_) );
OAI21X1 OAI21X1_3082 ( .A(_4763__bF_buf0), .B(_2240__bF_buf4), .C(_2258_), .Y(_588_) );
NAND2X1 NAND2X1_945 ( .A(cpuregs_25_[18]), .B(_2240__bF_buf3), .Y(_2259_) );
OAI21X1 OAI21X1_3083 ( .A(_4783__bF_buf0), .B(_2240__bF_buf2), .C(_2259_), .Y(_589_) );
NAND2X1 NAND2X1_946 ( .A(cpuregs_25_[19]), .B(_2240__bF_buf1), .Y(_2260_) );
OAI21X1 OAI21X1_3084 ( .A(_4793__bF_buf0), .B(_2240__bF_buf0), .C(_2260_), .Y(_590_) );
NAND2X1 NAND2X1_947 ( .A(cpuregs_25_[20]), .B(_2240__bF_buf7), .Y(_2261_) );
OAI21X1 OAI21X1_3085 ( .A(_4806__bF_buf0), .B(_2240__bF_buf6), .C(_2261_), .Y(_591_) );
NAND2X1 NAND2X1_948 ( .A(cpuregs_25_[21]), .B(_2240__bF_buf5), .Y(_2262_) );
OAI21X1 OAI21X1_3086 ( .A(_4816__bF_buf0), .B(_2240__bF_buf4), .C(_2262_), .Y(_592_) );
NAND2X1 NAND2X1_949 ( .A(cpuregs_25_[22]), .B(_2240__bF_buf3), .Y(_2263_) );
OAI21X1 OAI21X1_3087 ( .A(_4824__bF_buf0), .B(_2240__bF_buf2), .C(_2263_), .Y(_593_) );
NAND2X1 NAND2X1_950 ( .A(cpuregs_25_[23]), .B(_2240__bF_buf1), .Y(_2264_) );
OAI21X1 OAI21X1_3088 ( .A(_4833__bF_buf0), .B(_2240__bF_buf0), .C(_2264_), .Y(_594_) );
NAND2X1 NAND2X1_951 ( .A(cpuregs_25_[24]), .B(_2240__bF_buf7), .Y(_2265_) );
OAI21X1 OAI21X1_3089 ( .A(_4845__bF_buf0), .B(_2240__bF_buf6), .C(_2265_), .Y(_595_) );
NAND2X1 NAND2X1_952 ( .A(cpuregs_25_[25]), .B(_2240__bF_buf5), .Y(_2266_) );
OAI21X1 OAI21X1_3090 ( .A(_4854__bF_buf0), .B(_2240__bF_buf4), .C(_2266_), .Y(_596_) );
NAND2X1 NAND2X1_953 ( .A(cpuregs_25_[26]), .B(_2240__bF_buf3), .Y(_2267_) );
OAI21X1 OAI21X1_3091 ( .A(_4863__bF_buf0), .B(_2240__bF_buf2), .C(_2267_), .Y(_597_) );
NAND2X1 NAND2X1_954 ( .A(cpuregs_25_[27]), .B(_2240__bF_buf1), .Y(_2268_) );
OAI21X1 OAI21X1_3092 ( .A(_4871__bF_buf0), .B(_2240__bF_buf0), .C(_2268_), .Y(_598_) );
NAND2X1 NAND2X1_955 ( .A(cpuregs_25_[28]), .B(_2240__bF_buf7), .Y(_2269_) );
OAI21X1 OAI21X1_3093 ( .A(_4884__bF_buf0), .B(_2240__bF_buf6), .C(_2269_), .Y(_599_) );
NAND2X1 NAND2X1_956 ( .A(cpuregs_25_[29]), .B(_2240__bF_buf5), .Y(_2270_) );
OAI21X1 OAI21X1_3094 ( .A(_4893__bF_buf0), .B(_2240__bF_buf4), .C(_2270_), .Y(_600_) );
NAND2X1 NAND2X1_957 ( .A(cpuregs_25_[30]), .B(_2240__bF_buf3), .Y(_2271_) );
OAI21X1 OAI21X1_3095 ( .A(_4901__bF_buf0), .B(_2240__bF_buf2), .C(_2271_), .Y(_601_) );
NAND2X1 NAND2X1_958 ( .A(cpuregs_25_[31]), .B(_2240__bF_buf1), .Y(_2272_) );
OAI21X1 OAI21X1_3096 ( .A(_4910__bF_buf0), .B(_2240__bF_buf0), .C(_2272_), .Y(_602_) );
NOR2X1 NOR2X1_1222 ( .A(_2171__bF_buf5), .B(_5706__bF_buf5), .Y(_2273_) );
INVX1 INVX1_1177 ( .A(_2273_), .Y(_2274_) );
OAI21X1 OAI21X1_3097 ( .A(_5706__bF_buf4), .B(_2171__bF_buf4), .C(cpuregs_24_[0]), .Y(_2275_) );
OAI21X1 OAI21X1_3098 ( .A(_2274__bF_buf4), .B(_4925__bF_buf0), .C(_2275_), .Y(_603_) );
OAI21X1 OAI21X1_3099 ( .A(_5706__bF_buf3), .B(_2171__bF_buf3), .C(cpuregs_24_[1]), .Y(_2276_) );
OAI21X1 OAI21X1_3100 ( .A(_2274__bF_buf3), .B(_4933__bF_buf0), .C(_2276_), .Y(_604_) );
OAI21X1 OAI21X1_3101 ( .A(_5706__bF_buf2), .B(_2171__bF_buf2), .C(cpuregs_24_[2]), .Y(_2277_) );
OAI21X1 OAI21X1_3102 ( .A(_2274__bF_buf2), .B(_4940__bF_buf0), .C(_2277_), .Y(_605_) );
OAI21X1 OAI21X1_3103 ( .A(_5706__bF_buf1), .B(_2171__bF_buf1), .C(cpuregs_24_[3]), .Y(_2278_) );
OAI21X1 OAI21X1_3104 ( .A(_2274__bF_buf1), .B(_4948__bF_buf0), .C(_2278_), .Y(_606_) );
OAI21X1 OAI21X1_3105 ( .A(_5706__bF_buf0), .B(_2171__bF_buf0), .C(cpuregs_24_[4]), .Y(_2279_) );
OAI21X1 OAI21X1_3106 ( .A(_2274__bF_buf0), .B(_4955__bF_buf0), .C(_2279_), .Y(_607_) );
OAI21X1 OAI21X1_3107 ( .A(_5706__bF_buf11), .B(_2171__bF_buf8), .C(cpuregs_24_[5]), .Y(_2280_) );
OAI21X1 OAI21X1_3108 ( .A(_2274__bF_buf4), .B(_4654__bF_buf4), .C(_2280_), .Y(_608_) );
OAI21X1 OAI21X1_3109 ( .A(_5706__bF_buf10), .B(_2171__bF_buf7), .C(cpuregs_24_[6]), .Y(_2281_) );
OAI21X1 OAI21X1_3110 ( .A(_2274__bF_buf3), .B(_4664__bF_buf4), .C(_2281_), .Y(_609_) );
OAI21X1 OAI21X1_3111 ( .A(_5706__bF_buf9), .B(_2171__bF_buf6), .C(cpuregs_24_[7]), .Y(_2282_) );
OAI21X1 OAI21X1_3112 ( .A(_2274__bF_buf2), .B(_4677__bF_buf4), .C(_2282_), .Y(_610_) );
OAI21X1 OAI21X1_3113 ( .A(_5706__bF_buf8), .B(_2171__bF_buf5), .C(cpuregs_24_[8]), .Y(_2283_) );
OAI21X1 OAI21X1_3114 ( .A(_4685__bF_buf4), .B(_2274__bF_buf1), .C(_2283_), .Y(_611_) );
OAI21X1 OAI21X1_3115 ( .A(_5706__bF_buf7), .B(_2171__bF_buf4), .C(cpuregs_24_[9]), .Y(_2284_) );
OAI21X1 OAI21X1_3116 ( .A(_4696__bF_buf4), .B(_2274__bF_buf0), .C(_2284_), .Y(_612_) );
OAI21X1 OAI21X1_3117 ( .A(_5706__bF_buf6), .B(_2171__bF_buf3), .C(cpuregs_24_[10]), .Y(_2285_) );
OAI21X1 OAI21X1_3118 ( .A(_4703__bF_buf4), .B(_2274__bF_buf4), .C(_2285_), .Y(_613_) );
OAI21X1 OAI21X1_3119 ( .A(_5706__bF_buf5), .B(_2171__bF_buf2), .C(cpuregs_24_[11]), .Y(_2286_) );
OAI21X1 OAI21X1_3120 ( .A(_4713__bF_buf4), .B(_2274__bF_buf3), .C(_2286_), .Y(_614_) );
OAI21X1 OAI21X1_3121 ( .A(_5706__bF_buf4), .B(_2171__bF_buf1), .C(cpuregs_24_[12]), .Y(_2287_) );
OAI21X1 OAI21X1_3122 ( .A(_4722__bF_buf4), .B(_2274__bF_buf2), .C(_2287_), .Y(_615_) );
OAI21X1 OAI21X1_3123 ( .A(_5706__bF_buf3), .B(_2171__bF_buf0), .C(cpuregs_24_[13]), .Y(_2288_) );
OAI21X1 OAI21X1_3124 ( .A(_4731__bF_buf4), .B(_2274__bF_buf1), .C(_2288_), .Y(_616_) );
OAI21X1 OAI21X1_3125 ( .A(_5706__bF_buf2), .B(_2171__bF_buf8), .C(cpuregs_24_[14]), .Y(_2289_) );
OAI21X1 OAI21X1_3126 ( .A(_4740__bF_buf4), .B(_2274__bF_buf0), .C(_2289_), .Y(_617_) );
OAI21X1 OAI21X1_3127 ( .A(_5706__bF_buf1), .B(_2171__bF_buf7), .C(cpuregs_24_[15]), .Y(_2290_) );
OAI21X1 OAI21X1_3128 ( .A(_4747__bF_buf4), .B(_2274__bF_buf4), .C(_2290_), .Y(_618_) );
OAI21X1 OAI21X1_3129 ( .A(_5706__bF_buf0), .B(_2171__bF_buf6), .C(cpuregs_24_[16]), .Y(_2291_) );
OAI21X1 OAI21X1_3130 ( .A(_4755__bF_buf4), .B(_2274__bF_buf3), .C(_2291_), .Y(_619_) );
OAI21X1 OAI21X1_3131 ( .A(_5706__bF_buf11), .B(_2171__bF_buf5), .C(cpuregs_24_[17]), .Y(_2292_) );
OAI21X1 OAI21X1_3132 ( .A(_4763__bF_buf4), .B(_2274__bF_buf2), .C(_2292_), .Y(_620_) );
OAI21X1 OAI21X1_3133 ( .A(_5706__bF_buf10), .B(_2171__bF_buf4), .C(cpuregs_24_[18]), .Y(_2293_) );
OAI21X1 OAI21X1_3134 ( .A(_4783__bF_buf4), .B(_2274__bF_buf1), .C(_2293_), .Y(_621_) );
OAI21X1 OAI21X1_3135 ( .A(_5706__bF_buf9), .B(_2171__bF_buf3), .C(cpuregs_24_[19]), .Y(_2294_) );
OAI21X1 OAI21X1_3136 ( .A(_4793__bF_buf4), .B(_2274__bF_buf0), .C(_2294_), .Y(_622_) );
OAI21X1 OAI21X1_3137 ( .A(_5706__bF_buf8), .B(_2171__bF_buf2), .C(cpuregs_24_[20]), .Y(_2295_) );
OAI21X1 OAI21X1_3138 ( .A(_4806__bF_buf4), .B(_2274__bF_buf4), .C(_2295_), .Y(_623_) );
OAI21X1 OAI21X1_3139 ( .A(_5706__bF_buf7), .B(_2171__bF_buf1), .C(cpuregs_24_[21]), .Y(_2296_) );
OAI21X1 OAI21X1_3140 ( .A(_4816__bF_buf4), .B(_2274__bF_buf3), .C(_2296_), .Y(_624_) );
OAI21X1 OAI21X1_3141 ( .A(_5706__bF_buf6), .B(_2171__bF_buf0), .C(cpuregs_24_[22]), .Y(_2297_) );
OAI21X1 OAI21X1_3142 ( .A(_4824__bF_buf4), .B(_2274__bF_buf2), .C(_2297_), .Y(_625_) );
OAI21X1 OAI21X1_3143 ( .A(_5706__bF_buf5), .B(_2171__bF_buf8), .C(cpuregs_24_[23]), .Y(_2298_) );
OAI21X1 OAI21X1_3144 ( .A(_4833__bF_buf4), .B(_2274__bF_buf1), .C(_2298_), .Y(_626_) );
OAI21X1 OAI21X1_3145 ( .A(_5706__bF_buf4), .B(_2171__bF_buf7), .C(cpuregs_24_[24]), .Y(_2299_) );
OAI21X1 OAI21X1_3146 ( .A(_4845__bF_buf4), .B(_2274__bF_buf0), .C(_2299_), .Y(_627_) );
OAI21X1 OAI21X1_3147 ( .A(_5706__bF_buf3), .B(_2171__bF_buf6), .C(cpuregs_24_[25]), .Y(_2300_) );
OAI21X1 OAI21X1_3148 ( .A(_4854__bF_buf4), .B(_2274__bF_buf4), .C(_2300_), .Y(_628_) );
OAI21X1 OAI21X1_3149 ( .A(_5706__bF_buf2), .B(_2171__bF_buf5), .C(cpuregs_24_[26]), .Y(_2301_) );
OAI21X1 OAI21X1_3150 ( .A(_4863__bF_buf4), .B(_2274__bF_buf3), .C(_2301_), .Y(_629_) );
OAI21X1 OAI21X1_3151 ( .A(_5706__bF_buf1), .B(_2171__bF_buf4), .C(cpuregs_24_[27]), .Y(_2302_) );
OAI21X1 OAI21X1_3152 ( .A(_4871__bF_buf4), .B(_2274__bF_buf2), .C(_2302_), .Y(_630_) );
OAI21X1 OAI21X1_3153 ( .A(_5706__bF_buf0), .B(_2171__bF_buf3), .C(cpuregs_24_[28]), .Y(_2303_) );
OAI21X1 OAI21X1_3154 ( .A(_4884__bF_buf4), .B(_2274__bF_buf1), .C(_2303_), .Y(_631_) );
OAI21X1 OAI21X1_3155 ( .A(_5706__bF_buf11), .B(_2171__bF_buf2), .C(cpuregs_24_[29]), .Y(_2304_) );
OAI21X1 OAI21X1_3156 ( .A(_4893__bF_buf4), .B(_2274__bF_buf0), .C(_2304_), .Y(_632_) );
OAI21X1 OAI21X1_3157 ( .A(_5706__bF_buf10), .B(_2171__bF_buf1), .C(cpuregs_24_[30]), .Y(_2305_) );
OAI21X1 OAI21X1_3158 ( .A(_4901__bF_buf4), .B(_2274__bF_buf4), .C(_2305_), .Y(_633_) );
OAI21X1 OAI21X1_3159 ( .A(_5706__bF_buf9), .B(_2171__bF_buf0), .C(cpuregs_24_[31]), .Y(_2306_) );
OAI21X1 OAI21X1_3160 ( .A(_4910__bF_buf4), .B(_2274__bF_buf3), .C(_2306_), .Y(_634_) );
NOR2X1 NOR2X1_1223 ( .A(latched_rd_3_), .B(_5743_), .Y(_2307_) );
INVX1 INVX1_1178 ( .A(_2307_), .Y(_2308_) );
NOR2X1 NOR2X1_1224 ( .A(_4911_), .B(_2308_), .Y(_2309_) );
INVX1 INVX1_1179 ( .A(_2309_), .Y(_2310_) );
NOR2X1 NOR2X1_1225 ( .A(_2310__bF_buf7), .B(_4917__bF_buf10), .Y(_2311_) );
NOR2X1 NOR2X1_1226 ( .A(cpuregs_23_[0]), .B(_2311_), .Y(_2312_) );
AOI21X1 AOI21X1_913 ( .A(_4925__bF_buf4), .B(_2311_), .C(_2312_), .Y(_635_) );
NAND2X1 NAND2X1_959 ( .A(_4916_), .B(_2309_), .Y(_2313_) );
NOR2X1 NOR2X1_1227 ( .A(_2313__bF_buf3), .B(_4632__bF_buf0), .Y(_2314_) );
MUX2X1 MUX2X1_257 ( .A(_4933__bF_buf4), .B(_5480_), .S(_2314_), .Y(_636_) );
NOR2X1 NOR2X1_1228 ( .A(cpuregs_23_[2]), .B(_2311_), .Y(_2315_) );
AOI21X1 AOI21X1_914 ( .A(_4940__bF_buf4), .B(_2311_), .C(_2315_), .Y(_637_) );
MUX2X1 MUX2X1_258 ( .A(_4948__bF_buf4), .B(_5621_), .S(_2314_), .Y(_638_) );
NAND2X1 NAND2X1_960 ( .A(_2314_), .B(_5279_), .Y(_2316_) );
OAI21X1 OAI21X1_3161 ( .A(_5692_), .B(_2314_), .C(_2316_), .Y(_639_) );
NAND2X1 NAND2X1_961 ( .A(_2314_), .B(_4655_), .Y(_2317_) );
OAI21X1 OAI21X1_3162 ( .A(_5917_), .B(_2314_), .C(_2317_), .Y(_640_) );
NAND2X1 NAND2X1_962 ( .A(_2314_), .B(_4665_), .Y(_2318_) );
OAI21X1 OAI21X1_3163 ( .A(_5981_), .B(_2314_), .C(_2318_), .Y(_641_) );
INVX1 INVX1_1180 ( .A(_4677__bF_buf3), .Y(_2319_) );
NAND2X1 NAND2X1_963 ( .A(_2314_), .B(_2319_), .Y(_2320_) );
OAI21X1 OAI21X1_3164 ( .A(_6026_), .B(_2314_), .C(_2320_), .Y(_642_) );
NAND2X1 NAND2X1_964 ( .A(_2314_), .B(_4686_), .Y(_2321_) );
OAI21X1 OAI21X1_3165 ( .A(_6104_), .B(_2314_), .C(_2321_), .Y(_643_) );
NOR2X1 NOR2X1_1229 ( .A(cpuregs_23_[9]), .B(_2311_), .Y(_2322_) );
AOI21X1 AOI21X1_915 ( .A(_2311_), .B(_4696__bF_buf3), .C(_2322_), .Y(_644_) );
MUX2X1 MUX2X1_259 ( .A(_4703__bF_buf3), .B(_6210_), .S(_2311_), .Y(_645_) );
MUX2X1 MUX2X1_260 ( .A(_4713__bF_buf3), .B(_8397_), .S(_2311_), .Y(_646_) );
INVX1 INVX1_1181 ( .A(_2311_), .Y(_2323_) );
OAI21X1 OAI21X1_3166 ( .A(_4632__bF_buf8), .B(_2313__bF_buf2), .C(cpuregs_23_[12]), .Y(_2324_) );
OAI21X1 OAI21X1_3167 ( .A(_4722__bF_buf3), .B(_2323__bF_buf3), .C(_2324_), .Y(_647_) );
OAI21X1 OAI21X1_3168 ( .A(_4632__bF_buf7), .B(_2313__bF_buf1), .C(cpuregs_23_[13]), .Y(_2325_) );
OAI21X1 OAI21X1_3169 ( .A(_4731__bF_buf3), .B(_2323__bF_buf2), .C(_2325_), .Y(_648_) );
OAI21X1 OAI21X1_3170 ( .A(_4632__bF_buf6), .B(_2313__bF_buf0), .C(cpuregs_23_[14]), .Y(_2326_) );
OAI21X1 OAI21X1_3171 ( .A(_4740__bF_buf3), .B(_2323__bF_buf1), .C(_2326_), .Y(_649_) );
OAI21X1 OAI21X1_3172 ( .A(_4632__bF_buf5), .B(_2313__bF_buf3), .C(cpuregs_23_[15]), .Y(_2327_) );
OAI21X1 OAI21X1_3173 ( .A(_4747__bF_buf3), .B(_2323__bF_buf0), .C(_2327_), .Y(_650_) );
OAI21X1 OAI21X1_3174 ( .A(_4632__bF_buf4), .B(_2313__bF_buf2), .C(cpuregs_23_[16]), .Y(_2328_) );
OAI21X1 OAI21X1_3175 ( .A(_4755__bF_buf3), .B(_2323__bF_buf3), .C(_2328_), .Y(_651_) );
OAI21X1 OAI21X1_3176 ( .A(_4632__bF_buf3), .B(_2313__bF_buf1), .C(cpuregs_23_[17]), .Y(_2329_) );
OAI21X1 OAI21X1_3177 ( .A(_4763__bF_buf3), .B(_2323__bF_buf2), .C(_2329_), .Y(_652_) );
OAI21X1 OAI21X1_3178 ( .A(_4632__bF_buf2), .B(_2313__bF_buf0), .C(cpuregs_23_[18]), .Y(_2330_) );
OAI21X1 OAI21X1_3179 ( .A(_4783__bF_buf3), .B(_2323__bF_buf1), .C(_2330_), .Y(_653_) );
OAI21X1 OAI21X1_3180 ( .A(_4632__bF_buf1), .B(_2313__bF_buf3), .C(cpuregs_23_[19]), .Y(_2331_) );
OAI21X1 OAI21X1_3181 ( .A(_4793__bF_buf3), .B(_2323__bF_buf0), .C(_2331_), .Y(_654_) );
OAI21X1 OAI21X1_3182 ( .A(_4632__bF_buf0), .B(_2313__bF_buf2), .C(cpuregs_23_[20]), .Y(_2332_) );
OAI21X1 OAI21X1_3183 ( .A(_4806__bF_buf3), .B(_2323__bF_buf3), .C(_2332_), .Y(_655_) );
OAI21X1 OAI21X1_3184 ( .A(_4632__bF_buf8), .B(_2313__bF_buf1), .C(cpuregs_23_[21]), .Y(_2333_) );
OAI21X1 OAI21X1_3185 ( .A(_4816__bF_buf3), .B(_2323__bF_buf2), .C(_2333_), .Y(_656_) );
OAI21X1 OAI21X1_3186 ( .A(_4632__bF_buf7), .B(_2313__bF_buf0), .C(cpuregs_23_[22]), .Y(_2334_) );
OAI21X1 OAI21X1_3187 ( .A(_4824__bF_buf3), .B(_2323__bF_buf1), .C(_2334_), .Y(_657_) );
OAI21X1 OAI21X1_3188 ( .A(_4632__bF_buf6), .B(_2313__bF_buf3), .C(cpuregs_23_[23]), .Y(_2335_) );
OAI21X1 OAI21X1_3189 ( .A(_4833__bF_buf3), .B(_2323__bF_buf0), .C(_2335_), .Y(_658_) );
OAI21X1 OAI21X1_3190 ( .A(_4632__bF_buf5), .B(_2313__bF_buf2), .C(cpuregs_23_[24]), .Y(_2336_) );
OAI21X1 OAI21X1_3191 ( .A(_4845__bF_buf3), .B(_2323__bF_buf3), .C(_2336_), .Y(_659_) );
OAI21X1 OAI21X1_3192 ( .A(_4632__bF_buf4), .B(_2313__bF_buf1), .C(cpuregs_23_[25]), .Y(_2337_) );
OAI21X1 OAI21X1_3193 ( .A(_4854__bF_buf3), .B(_2323__bF_buf2), .C(_2337_), .Y(_660_) );
OAI21X1 OAI21X1_3194 ( .A(_4632__bF_buf3), .B(_2313__bF_buf0), .C(cpuregs_23_[26]), .Y(_2338_) );
OAI21X1 OAI21X1_3195 ( .A(_4863__bF_buf3), .B(_2323__bF_buf1), .C(_2338_), .Y(_661_) );
OAI21X1 OAI21X1_3196 ( .A(_4632__bF_buf2), .B(_2313__bF_buf3), .C(cpuregs_23_[27]), .Y(_2339_) );
OAI21X1 OAI21X1_3197 ( .A(_4871__bF_buf3), .B(_2323__bF_buf0), .C(_2339_), .Y(_662_) );
OAI21X1 OAI21X1_3198 ( .A(_4632__bF_buf1), .B(_2313__bF_buf2), .C(cpuregs_23_[28]), .Y(_2340_) );
OAI21X1 OAI21X1_3199 ( .A(_4884__bF_buf3), .B(_2323__bF_buf3), .C(_2340_), .Y(_663_) );
OAI21X1 OAI21X1_3200 ( .A(_4632__bF_buf0), .B(_2313__bF_buf1), .C(cpuregs_23_[29]), .Y(_2341_) );
OAI21X1 OAI21X1_3201 ( .A(_4893__bF_buf3), .B(_2323__bF_buf2), .C(_2341_), .Y(_664_) );
OAI21X1 OAI21X1_3202 ( .A(_4632__bF_buf8), .B(_2313__bF_buf0), .C(cpuregs_23_[30]), .Y(_2342_) );
OAI21X1 OAI21X1_3203 ( .A(_4901__bF_buf3), .B(_2323__bF_buf1), .C(_2342_), .Y(_665_) );
OAI21X1 OAI21X1_3204 ( .A(_4632__bF_buf7), .B(_2313__bF_buf3), .C(cpuregs_23_[31]), .Y(_2343_) );
OAI21X1 OAI21X1_3205 ( .A(_4910__bF_buf3), .B(_2323__bF_buf0), .C(_2343_), .Y(_666_) );
NOR2X1 NOR2X1_1230 ( .A(_2310__bF_buf6), .B(_5281__bF_buf8), .Y(_2344_) );
INVX1 INVX1_1182 ( .A(_2344_), .Y(_2345_) );
OAI21X1 OAI21X1_3206 ( .A(_5281__bF_buf7), .B(_2310__bF_buf5), .C(cpuregs_22_[0]), .Y(_2346_) );
OAI21X1 OAI21X1_3207 ( .A(_2345__bF_buf4), .B(_4925__bF_buf3), .C(_2346_), .Y(_667_) );
OAI21X1 OAI21X1_3208 ( .A(_5281__bF_buf6), .B(_2310__bF_buf4), .C(cpuregs_22_[1]), .Y(_2347_) );
OAI21X1 OAI21X1_3209 ( .A(_2345__bF_buf3), .B(_4933__bF_buf3), .C(_2347_), .Y(_668_) );
OAI21X1 OAI21X1_3210 ( .A(_5281__bF_buf5), .B(_2310__bF_buf3), .C(cpuregs_22_[2]), .Y(_2348_) );
OAI21X1 OAI21X1_3211 ( .A(_2345__bF_buf2), .B(_4940__bF_buf3), .C(_2348_), .Y(_669_) );
OAI21X1 OAI21X1_3212 ( .A(_5281__bF_buf4), .B(_2310__bF_buf2), .C(cpuregs_22_[3]), .Y(_2349_) );
OAI21X1 OAI21X1_3213 ( .A(_2345__bF_buf1), .B(_4948__bF_buf3), .C(_2349_), .Y(_670_) );
OAI21X1 OAI21X1_3214 ( .A(_5281__bF_buf3), .B(_2310__bF_buf1), .C(cpuregs_22_[4]), .Y(_2350_) );
OAI21X1 OAI21X1_3215 ( .A(_2345__bF_buf0), .B(_4955__bF_buf4), .C(_2350_), .Y(_671_) );
OAI21X1 OAI21X1_3216 ( .A(_5281__bF_buf2), .B(_2310__bF_buf0), .C(cpuregs_22_[5]), .Y(_2351_) );
OAI21X1 OAI21X1_3217 ( .A(_2345__bF_buf4), .B(_4654__bF_buf3), .C(_2351_), .Y(_672_) );
OAI21X1 OAI21X1_3218 ( .A(_5281__bF_buf1), .B(_2310__bF_buf7), .C(cpuregs_22_[6]), .Y(_2352_) );
OAI21X1 OAI21X1_3219 ( .A(_4664__bF_buf3), .B(_2345__bF_buf3), .C(_2352_), .Y(_673_) );
OAI21X1 OAI21X1_3220 ( .A(_5281__bF_buf0), .B(_2310__bF_buf6), .C(cpuregs_22_[7]), .Y(_2353_) );
OAI21X1 OAI21X1_3221 ( .A(_4677__bF_buf2), .B(_2345__bF_buf2), .C(_2353_), .Y(_674_) );
OAI21X1 OAI21X1_3222 ( .A(_5281__bF_buf10), .B(_2310__bF_buf5), .C(cpuregs_22_[8]), .Y(_2354_) );
OAI21X1 OAI21X1_3223 ( .A(_4685__bF_buf3), .B(_2345__bF_buf1), .C(_2354_), .Y(_675_) );
OAI21X1 OAI21X1_3224 ( .A(_5281__bF_buf9), .B(_2310__bF_buf4), .C(cpuregs_22_[9]), .Y(_2355_) );
OAI21X1 OAI21X1_3225 ( .A(_4696__bF_buf2), .B(_2345__bF_buf0), .C(_2355_), .Y(_676_) );
OAI21X1 OAI21X1_3226 ( .A(_5281__bF_buf8), .B(_2310__bF_buf3), .C(cpuregs_22_[10]), .Y(_2356_) );
OAI21X1 OAI21X1_3227 ( .A(_4703__bF_buf2), .B(_2345__bF_buf4), .C(_2356_), .Y(_677_) );
OAI21X1 OAI21X1_3228 ( .A(_5281__bF_buf7), .B(_2310__bF_buf2), .C(cpuregs_22_[11]), .Y(_2357_) );
OAI21X1 OAI21X1_3229 ( .A(_4713__bF_buf2), .B(_2345__bF_buf3), .C(_2357_), .Y(_678_) );
OAI21X1 OAI21X1_3230 ( .A(_5281__bF_buf6), .B(_2310__bF_buf1), .C(cpuregs_22_[12]), .Y(_2358_) );
OAI21X1 OAI21X1_3231 ( .A(_4722__bF_buf2), .B(_2345__bF_buf2), .C(_2358_), .Y(_679_) );
OAI21X1 OAI21X1_3232 ( .A(_5281__bF_buf5), .B(_2310__bF_buf0), .C(cpuregs_22_[13]), .Y(_2359_) );
OAI21X1 OAI21X1_3233 ( .A(_4731__bF_buf2), .B(_2345__bF_buf1), .C(_2359_), .Y(_680_) );
OAI21X1 OAI21X1_3234 ( .A(_5281__bF_buf4), .B(_2310__bF_buf7), .C(cpuregs_22_[14]), .Y(_2360_) );
OAI21X1 OAI21X1_3235 ( .A(_4740__bF_buf2), .B(_2345__bF_buf0), .C(_2360_), .Y(_681_) );
OAI21X1 OAI21X1_3236 ( .A(_5281__bF_buf3), .B(_2310__bF_buf6), .C(cpuregs_22_[15]), .Y(_2361_) );
OAI21X1 OAI21X1_3237 ( .A(_4747__bF_buf2), .B(_2345__bF_buf4), .C(_2361_), .Y(_682_) );
OAI21X1 OAI21X1_3238 ( .A(_5281__bF_buf2), .B(_2310__bF_buf5), .C(cpuregs_22_[16]), .Y(_2362_) );
OAI21X1 OAI21X1_3239 ( .A(_4755__bF_buf2), .B(_2345__bF_buf3), .C(_2362_), .Y(_683_) );
OAI21X1 OAI21X1_3240 ( .A(_5281__bF_buf1), .B(_2310__bF_buf4), .C(cpuregs_22_[17]), .Y(_2363_) );
OAI21X1 OAI21X1_3241 ( .A(_4763__bF_buf2), .B(_2345__bF_buf2), .C(_2363_), .Y(_684_) );
OAI21X1 OAI21X1_3242 ( .A(_5281__bF_buf0), .B(_2310__bF_buf3), .C(cpuregs_22_[18]), .Y(_2364_) );
OAI21X1 OAI21X1_3243 ( .A(_4783__bF_buf2), .B(_2345__bF_buf1), .C(_2364_), .Y(_685_) );
OAI21X1 OAI21X1_3244 ( .A(_5281__bF_buf10), .B(_2310__bF_buf2), .C(cpuregs_22_[19]), .Y(_2365_) );
OAI21X1 OAI21X1_3245 ( .A(_4793__bF_buf2), .B(_2345__bF_buf0), .C(_2365_), .Y(_686_) );
OAI21X1 OAI21X1_3246 ( .A(_5281__bF_buf9), .B(_2310__bF_buf1), .C(cpuregs_22_[20]), .Y(_2366_) );
OAI21X1 OAI21X1_3247 ( .A(_4806__bF_buf2), .B(_2345__bF_buf4), .C(_2366_), .Y(_687_) );
OAI21X1 OAI21X1_3248 ( .A(_5281__bF_buf8), .B(_2310__bF_buf0), .C(cpuregs_22_[21]), .Y(_2367_) );
OAI21X1 OAI21X1_3249 ( .A(_4816__bF_buf2), .B(_2345__bF_buf3), .C(_2367_), .Y(_688_) );
OAI21X1 OAI21X1_3250 ( .A(_5281__bF_buf7), .B(_2310__bF_buf7), .C(cpuregs_22_[22]), .Y(_2368_) );
OAI21X1 OAI21X1_3251 ( .A(_4824__bF_buf2), .B(_2345__bF_buf2), .C(_2368_), .Y(_689_) );
OAI21X1 OAI21X1_3252 ( .A(_5281__bF_buf6), .B(_2310__bF_buf6), .C(cpuregs_22_[23]), .Y(_2369_) );
OAI21X1 OAI21X1_3253 ( .A(_4833__bF_buf2), .B(_2345__bF_buf1), .C(_2369_), .Y(_690_) );
OAI21X1 OAI21X1_3254 ( .A(_5281__bF_buf5), .B(_2310__bF_buf5), .C(cpuregs_22_[24]), .Y(_2370_) );
OAI21X1 OAI21X1_3255 ( .A(_4845__bF_buf2), .B(_2345__bF_buf0), .C(_2370_), .Y(_691_) );
OAI21X1 OAI21X1_3256 ( .A(_5281__bF_buf4), .B(_2310__bF_buf4), .C(cpuregs_22_[25]), .Y(_2371_) );
OAI21X1 OAI21X1_3257 ( .A(_4854__bF_buf2), .B(_2345__bF_buf4), .C(_2371_), .Y(_692_) );
OAI21X1 OAI21X1_3258 ( .A(_5281__bF_buf3), .B(_2310__bF_buf3), .C(cpuregs_22_[26]), .Y(_2372_) );
OAI21X1 OAI21X1_3259 ( .A(_4863__bF_buf2), .B(_2345__bF_buf3), .C(_2372_), .Y(_693_) );
OAI21X1 OAI21X1_3260 ( .A(_5281__bF_buf2), .B(_2310__bF_buf2), .C(cpuregs_22_[27]), .Y(_2373_) );
OAI21X1 OAI21X1_3261 ( .A(_4871__bF_buf2), .B(_2345__bF_buf2), .C(_2373_), .Y(_694_) );
OAI21X1 OAI21X1_3262 ( .A(_5281__bF_buf1), .B(_2310__bF_buf1), .C(cpuregs_22_[28]), .Y(_2374_) );
OAI21X1 OAI21X1_3263 ( .A(_4884__bF_buf2), .B(_2345__bF_buf1), .C(_2374_), .Y(_695_) );
OAI21X1 OAI21X1_3264 ( .A(_5281__bF_buf0), .B(_2310__bF_buf0), .C(cpuregs_22_[29]), .Y(_2375_) );
OAI21X1 OAI21X1_3265 ( .A(_4893__bF_buf2), .B(_2345__bF_buf0), .C(_2375_), .Y(_696_) );
OAI21X1 OAI21X1_3266 ( .A(_5281__bF_buf10), .B(_2310__bF_buf7), .C(cpuregs_22_[30]), .Y(_2376_) );
OAI21X1 OAI21X1_3267 ( .A(_4901__bF_buf2), .B(_2345__bF_buf4), .C(_2376_), .Y(_697_) );
OAI21X1 OAI21X1_3268 ( .A(_5281__bF_buf9), .B(_2310__bF_buf6), .C(cpuregs_22_[31]), .Y(_2377_) );
OAI21X1 OAI21X1_3269 ( .A(_4910__bF_buf2), .B(_2345__bF_buf3), .C(_2377_), .Y(_698_) );
NAND2X1 NAND2X1_965 ( .A(_2309_), .B(_5313_), .Y(_2378_) );
NAND2X1 NAND2X1_966 ( .A(cpuregs_21_[0]), .B(_2378__bF_buf7), .Y(_2379_) );
OAI21X1 OAI21X1_3270 ( .A(_4925__bF_buf2), .B(_2378__bF_buf6), .C(_2379_), .Y(_699_) );
NAND2X1 NAND2X1_967 ( .A(cpuregs_21_[1]), .B(_2378__bF_buf5), .Y(_2380_) );
OAI21X1 OAI21X1_3271 ( .A(_4933__bF_buf2), .B(_2378__bF_buf4), .C(_2380_), .Y(_700_) );
NAND2X1 NAND2X1_968 ( .A(cpuregs_21_[2]), .B(_2378__bF_buf3), .Y(_2381_) );
OAI21X1 OAI21X1_3272 ( .A(_4940__bF_buf2), .B(_2378__bF_buf2), .C(_2381_), .Y(_701_) );
NAND2X1 NAND2X1_969 ( .A(cpuregs_21_[3]), .B(_2378__bF_buf1), .Y(_2382_) );
OAI21X1 OAI21X1_3273 ( .A(_4948__bF_buf2), .B(_2378__bF_buf0), .C(_2382_), .Y(_702_) );
NAND2X1 NAND2X1_970 ( .A(cpuregs_21_[4]), .B(_2378__bF_buf7), .Y(_2383_) );
OAI21X1 OAI21X1_3274 ( .A(_4955__bF_buf3), .B(_2378__bF_buf6), .C(_2383_), .Y(_703_) );
NAND2X1 NAND2X1_971 ( .A(cpuregs_21_[5]), .B(_2378__bF_buf5), .Y(_2384_) );
OAI21X1 OAI21X1_3275 ( .A(_4654__bF_buf2), .B(_2378__bF_buf4), .C(_2384_), .Y(_704_) );
NAND2X1 NAND2X1_972 ( .A(cpuregs_21_[6]), .B(_2378__bF_buf3), .Y(_2385_) );
OAI21X1 OAI21X1_3276 ( .A(_4664__bF_buf2), .B(_2378__bF_buf2), .C(_2385_), .Y(_705_) );
NAND2X1 NAND2X1_973 ( .A(cpuregs_21_[7]), .B(_2378__bF_buf1), .Y(_2386_) );
OAI21X1 OAI21X1_3277 ( .A(_4677__bF_buf1), .B(_2378__bF_buf0), .C(_2386_), .Y(_706_) );
NAND2X1 NAND2X1_974 ( .A(cpuregs_21_[8]), .B(_2378__bF_buf7), .Y(_2387_) );
OAI21X1 OAI21X1_3278 ( .A(_4685__bF_buf2), .B(_2378__bF_buf6), .C(_2387_), .Y(_707_) );
NAND2X1 NAND2X1_975 ( .A(cpuregs_21_[9]), .B(_2378__bF_buf5), .Y(_2388_) );
OAI21X1 OAI21X1_3279 ( .A(_4696__bF_buf1), .B(_2378__bF_buf4), .C(_2388_), .Y(_708_) );
NAND2X1 NAND2X1_976 ( .A(cpuregs_21_[10]), .B(_2378__bF_buf3), .Y(_2389_) );
OAI21X1 OAI21X1_3280 ( .A(_4703__bF_buf1), .B(_2378__bF_buf2), .C(_2389_), .Y(_709_) );
NAND2X1 NAND2X1_977 ( .A(cpuregs_21_[11]), .B(_2378__bF_buf1), .Y(_2390_) );
OAI21X1 OAI21X1_3281 ( .A(_4713__bF_buf1), .B(_2378__bF_buf0), .C(_2390_), .Y(_710_) );
NAND2X1 NAND2X1_978 ( .A(cpuregs_21_[12]), .B(_2378__bF_buf7), .Y(_2391_) );
OAI21X1 OAI21X1_3282 ( .A(_4722__bF_buf1), .B(_2378__bF_buf6), .C(_2391_), .Y(_711_) );
NAND2X1 NAND2X1_979 ( .A(cpuregs_21_[13]), .B(_2378__bF_buf5), .Y(_2392_) );
OAI21X1 OAI21X1_3283 ( .A(_4731__bF_buf1), .B(_2378__bF_buf4), .C(_2392_), .Y(_712_) );
NAND2X1 NAND2X1_980 ( .A(cpuregs_21_[14]), .B(_2378__bF_buf3), .Y(_2393_) );
OAI21X1 OAI21X1_3284 ( .A(_4740__bF_buf1), .B(_2378__bF_buf2), .C(_2393_), .Y(_713_) );
NAND2X1 NAND2X1_981 ( .A(cpuregs_21_[15]), .B(_2378__bF_buf1), .Y(_2394_) );
OAI21X1 OAI21X1_3285 ( .A(_4747__bF_buf1), .B(_2378__bF_buf0), .C(_2394_), .Y(_714_) );
NAND2X1 NAND2X1_982 ( .A(cpuregs_21_[16]), .B(_2378__bF_buf7), .Y(_2395_) );
OAI21X1 OAI21X1_3286 ( .A(_4755__bF_buf1), .B(_2378__bF_buf6), .C(_2395_), .Y(_715_) );
NAND2X1 NAND2X1_983 ( .A(cpuregs_21_[17]), .B(_2378__bF_buf5), .Y(_2396_) );
OAI21X1 OAI21X1_3287 ( .A(_4763__bF_buf1), .B(_2378__bF_buf4), .C(_2396_), .Y(_716_) );
NAND2X1 NAND2X1_984 ( .A(cpuregs_21_[18]), .B(_2378__bF_buf3), .Y(_2397_) );
OAI21X1 OAI21X1_3288 ( .A(_4783__bF_buf1), .B(_2378__bF_buf2), .C(_2397_), .Y(_717_) );
NAND2X1 NAND2X1_985 ( .A(cpuregs_21_[19]), .B(_2378__bF_buf1), .Y(_2398_) );
OAI21X1 OAI21X1_3289 ( .A(_4793__bF_buf1), .B(_2378__bF_buf0), .C(_2398_), .Y(_718_) );
NAND2X1 NAND2X1_986 ( .A(cpuregs_21_[20]), .B(_2378__bF_buf7), .Y(_2399_) );
OAI21X1 OAI21X1_3290 ( .A(_4806__bF_buf1), .B(_2378__bF_buf6), .C(_2399_), .Y(_719_) );
NAND2X1 NAND2X1_987 ( .A(cpuregs_21_[21]), .B(_2378__bF_buf5), .Y(_2400_) );
OAI21X1 OAI21X1_3291 ( .A(_4816__bF_buf1), .B(_2378__bF_buf4), .C(_2400_), .Y(_720_) );
NAND2X1 NAND2X1_988 ( .A(cpuregs_21_[22]), .B(_2378__bF_buf3), .Y(_2401_) );
OAI21X1 OAI21X1_3292 ( .A(_4824__bF_buf1), .B(_2378__bF_buf2), .C(_2401_), .Y(_721_) );
NAND2X1 NAND2X1_989 ( .A(cpuregs_21_[23]), .B(_2378__bF_buf1), .Y(_2402_) );
OAI21X1 OAI21X1_3293 ( .A(_4833__bF_buf1), .B(_2378__bF_buf0), .C(_2402_), .Y(_722_) );
NAND2X1 NAND2X1_990 ( .A(cpuregs_21_[24]), .B(_2378__bF_buf7), .Y(_2403_) );
OAI21X1 OAI21X1_3294 ( .A(_4845__bF_buf1), .B(_2378__bF_buf6), .C(_2403_), .Y(_723_) );
NAND2X1 NAND2X1_991 ( .A(cpuregs_21_[25]), .B(_2378__bF_buf5), .Y(_2404_) );
OAI21X1 OAI21X1_3295 ( .A(_4854__bF_buf1), .B(_2378__bF_buf4), .C(_2404_), .Y(_724_) );
NAND2X1 NAND2X1_992 ( .A(cpuregs_21_[26]), .B(_2378__bF_buf3), .Y(_2405_) );
OAI21X1 OAI21X1_3296 ( .A(_4863__bF_buf1), .B(_2378__bF_buf2), .C(_2405_), .Y(_725_) );
NAND2X1 NAND2X1_993 ( .A(cpuregs_21_[27]), .B(_2378__bF_buf1), .Y(_2406_) );
OAI21X1 OAI21X1_3297 ( .A(_4871__bF_buf1), .B(_2378__bF_buf0), .C(_2406_), .Y(_726_) );
NAND2X1 NAND2X1_994 ( .A(cpuregs_21_[28]), .B(_2378__bF_buf7), .Y(_2407_) );
OAI21X1 OAI21X1_3298 ( .A(_4884__bF_buf1), .B(_2378__bF_buf6), .C(_2407_), .Y(_727_) );
NAND2X1 NAND2X1_995 ( .A(cpuregs_21_[29]), .B(_2378__bF_buf5), .Y(_2408_) );
OAI21X1 OAI21X1_3299 ( .A(_4893__bF_buf1), .B(_2378__bF_buf4), .C(_2408_), .Y(_728_) );
NAND2X1 NAND2X1_996 ( .A(cpuregs_21_[30]), .B(_2378__bF_buf3), .Y(_2409_) );
OAI21X1 OAI21X1_3300 ( .A(_4901__bF_buf1), .B(_2378__bF_buf2), .C(_2409_), .Y(_729_) );
NAND2X1 NAND2X1_997 ( .A(cpuregs_21_[31]), .B(_2378__bF_buf1), .Y(_2410_) );
OAI21X1 OAI21X1_3301 ( .A(_4910__bF_buf1), .B(_2378__bF_buf0), .C(_2410_), .Y(_730_) );
NOR2X1 NOR2X1_1231 ( .A(_4923_), .B(_7620_), .Y(_2411_) );
OAI21X1 OAI21X1_3302 ( .A(reg_pc_0_), .B(decoded_imm_0_), .C(cpu_state_3_bF_buf2_), .Y(_2412_) );
NOR2X1 NOR2X1_1232 ( .A(_10734__1_), .B(_4491_), .Y(_2413_) );
NOR2X1 NOR2X1_1233 ( .A(_4490_), .B(_4491_), .Y(_2414_) );
AOI22X1 AOI22X1_129 ( .A(_2413_), .B(mem_rdata[8]), .C(mem_rdata[24]), .D(_2414_), .Y(_2415_) );
NOR2X1 NOR2X1_1234 ( .A(_1817__bF_buf0), .B(_2415_), .Y(_2416_) );
INVX1 INVX1_1183 ( .A(_10730__0_), .Y(_2417_) );
NAND2X1 NAND2X1_998 ( .A(mem_rdata[16]), .B(_1809_), .Y(_2418_) );
OAI21X1 OAI21X1_3303 ( .A(_2417_), .B(_1549_), .C(_2418_), .Y(_2419_) );
OR2X2 OR2X2_41 ( .A(_2419_), .B(_2416_), .Y(_2420_) );
INVX1 INVX1_1184 ( .A(_4531__bF_buf3), .Y(_2421_) );
INVX1 INVX1_1185 ( .A(count_instr_0_), .Y(_2422_) );
AOI22X1 AOI22X1_130 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_0_), .C(instr_rdcycleh_bF_buf1), .D(count_cycle_32_), .Y(_2423_) );
OAI21X1 OAI21X1_3304 ( .A(_4529_), .B(_2422_), .C(_2423_), .Y(_2424_) );
AOI21X1 AOI21X1_916 ( .A(count_instr_32_), .B(_2421_), .C(_2424_), .Y(_2425_) );
OAI22X1 OAI22X1_272 ( .A(_4575__bF_buf1), .B(_4491_), .C(_2425_), .D(_4538__bF_buf0), .Y(_2426_) );
AOI21X1 AOI21X1_917 ( .A(_4447__bF_buf1), .B(_2420_), .C(_2426_), .Y(_2427_) );
OAI21X1 OAI21X1_3305 ( .A(_2411_), .B(_2412_), .C(_2427_), .Y(_83__0_) );
NOR2X1 NOR2X1_1235 ( .A(_1541_), .B(_1810_), .Y(_2428_) );
AOI22X1 AOI22X1_131 ( .A(_2413_), .B(mem_rdata[9]), .C(mem_rdata[25]), .D(_2414_), .Y(_2429_) );
OAI22X1 OAI22X1_273 ( .A(_1817__bF_buf3), .B(_2429_), .C(_2417_), .D(_1551_), .Y(_2430_) );
OAI21X1 OAI21X1_3306 ( .A(_2430_), .B(_2428_), .C(_4447__bF_buf0), .Y(_2431_) );
INVX1 INVX1_1186 ( .A(_2411_), .Y(_2432_) );
XNOR2X1 XNOR2X1_50 ( .A(reg_pc_1_), .B(decoded_imm_1_), .Y(_2433_) );
AOI21X1 AOI21X1_918 ( .A(_2433_), .B(_2432_), .C(_4555_), .Y(_2434_) );
OAI21X1 OAI21X1_3307 ( .A(_2432_), .B(_2433_), .C(_2434_), .Y(_2435_) );
NAND2X1 NAND2X1_999 ( .A(instr_rdinstr_bF_buf3), .B(count_instr_1_), .Y(_2436_) );
AOI22X1 AOI22X1_132 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_1_), .C(instr_rdcycleh_bF_buf0), .D(count_cycle_33_), .Y(_2437_) );
NAND3X1 NAND3X1_94 ( .A(_2436_), .B(_2437_), .C(_4531__bF_buf2), .Y(_2438_) );
OAI21X1 OAI21X1_3308 ( .A(count_instr_33_), .B(_4531__bF_buf1), .C(_2438_), .Y(_2439_) );
NOR2X1 NOR2X1_1236 ( .A(_4538__bF_buf4), .B(_2439_), .Y(_2440_) );
AOI21X1 AOI21X1_919 ( .A(cpu_state_4_), .B(_10734__1_), .C(_2440_), .Y(_2441_) );
NAND3X1 NAND3X1_95 ( .A(_2435_), .B(_2441_), .C(_2431_), .Y(_83__1_) );
AOI22X1 AOI22X1_133 ( .A(_2413_), .B(mem_rdata[10]), .C(mem_rdata[26]), .D(_2414_), .Y(_2442_) );
NOR2X1 NOR2X1_1237 ( .A(_1817__bF_buf2), .B(_2442_), .Y(_2443_) );
OAI22X1 OAI22X1_274 ( .A(_1544_), .B(_1810_), .C(_2417_), .D(_4549_), .Y(_2444_) );
OAI21X1 OAI21X1_3309 ( .A(_2444_), .B(_2443_), .C(_4447__bF_buf3), .Y(_2445_) );
NOR2X1 NOR2X1_1238 ( .A(_2433_), .B(_2432_), .Y(_2446_) );
AOI21X1 AOI21X1_920 ( .A(reg_pc_1_), .B(decoded_imm_1_), .C(_2446_), .Y(_2447_) );
NAND2X1 NAND2X1_1000 ( .A(_4644_), .B(_7766_), .Y(_2448_) );
NAND2X1 NAND2X1_1001 ( .A(reg_pc_2_), .B(decoded_imm_2_), .Y(_2449_) );
NAND2X1 NAND2X1_1002 ( .A(_2449_), .B(_2448_), .Y(_2450_) );
OAI21X1 OAI21X1_3310 ( .A(_2447_), .B(_2450_), .C(cpu_state_3_bF_buf1_), .Y(_2451_) );
AOI21X1 AOI21X1_921 ( .A(_2447_), .B(_2450_), .C(_2451_), .Y(_2452_) );
INVX1 INVX1_1187 ( .A(count_cycle_34_), .Y(_2453_) );
AOI22X1 AOI22X1_134 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_2_), .C(instr_rdinstr_bF_buf2), .D(count_instr_2_), .Y(_2454_) );
OAI21X1 OAI21X1_3311 ( .A(_1735_), .B(_2453_), .C(_2454_), .Y(_2455_) );
AOI21X1 AOI21X1_922 ( .A(count_instr_34_), .B(_2421_), .C(_2455_), .Y(_2456_) );
OAI22X1 OAI22X1_275 ( .A(_4575__bF_buf0), .B(_5148_), .C(_2456_), .D(_4538__bF_buf3), .Y(_2457_) );
NOR2X1 NOR2X1_1239 ( .A(_2457_), .B(_2452_), .Y(_2458_) );
NAND2X1 NAND2X1_1003 ( .A(_2445_), .B(_2458_), .Y(_83__2_) );
OAI21X1 OAI21X1_3312 ( .A(_2447_), .B(_2450_), .C(_2449_), .Y(_2459_) );
NOR2X1 NOR2X1_1240 ( .A(reg_pc_3_), .B(decoded_imm_3_), .Y(_2460_) );
NOR2X1 NOR2X1_1241 ( .A(_7786_), .B(_7850_), .Y(_2461_) );
NOR2X1 NOR2X1_1242 ( .A(_2460_), .B(_2461_), .Y(_2462_) );
AND2X2 AND2X2_201 ( .A(_2459_), .B(_2462_), .Y(_2463_) );
OAI21X1 OAI21X1_3313 ( .A(_2459_), .B(_2462_), .C(cpu_state_3_bF_buf0_), .Y(_2464_) );
NOR2X1 NOR2X1_1243 ( .A(_10734__1_), .B(_10734__0_), .Y(_2465_) );
OAI21X1 OAI21X1_3314 ( .A(_1798_), .B(_2465_), .C(mem_rdata[3]), .Y(_2466_) );
INVX1 INVX1_1188 ( .A(_2413_), .Y(_2467_) );
NAND2X1 NAND2X1_1004 ( .A(mem_rdata[27]), .B(_2414_), .Y(_2468_) );
OAI21X1 OAI21X1_3315 ( .A(_2467_), .B(_1702_), .C(_2468_), .Y(_2469_) );
AOI22X1 AOI22X1_135 ( .A(mem_rdata[19]), .B(_1809_), .C(_2469_), .D(_1816_), .Y(_2470_) );
NAND2X1 NAND2X1_1005 ( .A(_2466_), .B(_2470_), .Y(_2471_) );
NOR2X1 NOR2X1_1244 ( .A(_1362_), .B(_4531__bF_buf0), .Y(_2472_) );
NAND2X1 NAND2X1_1006 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_3_), .Y(_2473_) );
NAND2X1 NAND2X1_1007 ( .A(instr_rdinstr_bF_buf1), .B(count_instr_3_), .Y(_2474_) );
NAND2X1 NAND2X1_1008 ( .A(instr_rdcycleh_bF_buf3), .B(count_cycle_35_), .Y(_2475_) );
NAND3X1 NAND3X1_96 ( .A(_2473_), .B(_2474_), .C(_2475_), .Y(_2476_) );
OAI21X1 OAI21X1_3316 ( .A(_2472_), .B(_2476_), .C(cpu_state_2_bF_buf2_), .Y(_2477_) );
OAI21X1 OAI21X1_3317 ( .A(_4575__bF_buf4), .B(_5130_), .C(_2477_), .Y(_2478_) );
AOI21X1 AOI21X1_923 ( .A(_4447__bF_buf2), .B(_2471_), .C(_2478_), .Y(_2479_) );
OAI21X1 OAI21X1_3318 ( .A(_2463_), .B(_2464_), .C(_2479_), .Y(_83__3_) );
NAND2X1 NAND2X1_1009 ( .A(_4642_), .B(_7914_), .Y(_2480_) );
NOR2X1 NOR2X1_1245 ( .A(_4642_), .B(_7914_), .Y(_2481_) );
INVX1 INVX1_1189 ( .A(_2481_), .Y(_2482_) );
NAND2X1 NAND2X1_1010 ( .A(_2480_), .B(_2482_), .Y(_2483_) );
INVX1 INVX1_1190 ( .A(_2460_), .Y(_2484_) );
AOI21X1 AOI21X1_924 ( .A(_2484_), .B(_2459_), .C(_2461_), .Y(_2485_) );
XNOR2X1 XNOR2X1_51 ( .A(_2485_), .B(_2483_), .Y(_2486_) );
AOI22X1 AOI22X1_136 ( .A(_2413_), .B(mem_rdata[12]), .C(mem_rdata[28]), .D(_2414_), .Y(_2487_) );
AOI22X1 AOI22X1_137 ( .A(mem_rdata[20]), .B(_1809_), .C(_10730__0_), .D(mem_rdata[4]), .Y(_2488_) );
OAI21X1 OAI21X1_3319 ( .A(_2487_), .B(_1817__bF_buf1), .C(_2488_), .Y(_2489_) );
NOR2X1 NOR2X1_1246 ( .A(_1368_), .B(_4531__bF_buf4), .Y(_2490_) );
NAND2X1 NAND2X1_1011 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_4_), .Y(_2491_) );
NAND2X1 NAND2X1_1012 ( .A(instr_rdinstr_bF_buf0), .B(count_instr_4_), .Y(_2492_) );
NAND2X1 NAND2X1_1013 ( .A(instr_rdcycleh_bF_buf2), .B(count_cycle_36_), .Y(_2493_) );
NAND3X1 NAND3X1_97 ( .A(_2491_), .B(_2492_), .C(_2493_), .Y(_2494_) );
OAI21X1 OAI21X1_3320 ( .A(_2490_), .B(_2494_), .C(cpu_state_2_bF_buf1_), .Y(_2495_) );
OAI21X1 OAI21X1_3321 ( .A(_4575__bF_buf3), .B(_5180_), .C(_2495_), .Y(_2496_) );
AOI21X1 AOI21X1_925 ( .A(_4447__bF_buf1), .B(_2489_), .C(_2496_), .Y(_2497_) );
OAI21X1 OAI21X1_3322 ( .A(_2486_), .B(_4555_), .C(_2497_), .Y(_83__4_) );
NAND2X1 NAND2X1_1014 ( .A(mem_rdata[29]), .B(_2414_), .Y(_2498_) );
OAI21X1 OAI21X1_3323 ( .A(_2467_), .B(_4615_), .C(_2498_), .Y(_2499_) );
INVX1 INVX1_1191 ( .A(mem_rdata[21]), .Y(_2500_) );
OAI21X1 OAI21X1_3324 ( .A(_1798_), .B(_2465_), .C(mem_rdata[5]), .Y(_2501_) );
OAI21X1 OAI21X1_3325 ( .A(_1810_), .B(_2500_), .C(_2501_), .Y(_2502_) );
AOI21X1 AOI21X1_926 ( .A(_1816_), .B(_2499_), .C(_2502_), .Y(_2503_) );
XNOR2X1 XNOR2X1_52 ( .A(reg_pc_5_), .B(decoded_imm_5_), .Y(_2504_) );
OAI21X1 OAI21X1_3326 ( .A(_2485_), .B(_2483_), .C(_2482_), .Y(_2505_) );
XNOR2X1 XNOR2X1_53 ( .A(_2505_), .B(_2504_), .Y(_2506_) );
NOR2X1 NOR2X1_1247 ( .A(_1372_), .B(_4531__bF_buf3), .Y(_2507_) );
INVX1 INVX1_1192 ( .A(count_cycle_37_), .Y(_2508_) );
AOI22X1 AOI22X1_138 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_5_), .C(instr_rdinstr_bF_buf4), .D(count_instr_5_), .Y(_2509_) );
OAI21X1 OAI21X1_3327 ( .A(_1735_), .B(_2508_), .C(_2509_), .Y(_2510_) );
OAI21X1 OAI21X1_3328 ( .A(_2507_), .B(_2510_), .C(cpu_state_2_bF_buf0_), .Y(_2511_) );
OAI21X1 OAI21X1_3329 ( .A(_4575__bF_buf2), .B(_5179_), .C(_2511_), .Y(_2512_) );
AOI21X1 AOI21X1_927 ( .A(cpu_state_3_bF_buf4_), .B(_2506_), .C(_2512_), .Y(_2513_) );
OAI21X1 OAI21X1_3330 ( .A(_4448_), .B(_2503_), .C(_2513_), .Y(_83__5_) );
NOR2X1 NOR2X1_1248 ( .A(_2504_), .B(_2483_), .Y(_2514_) );
INVX1 INVX1_1193 ( .A(_2514_), .Y(_2515_) );
NOR2X1 NOR2X1_1249 ( .A(_2504_), .B(_2482_), .Y(_2516_) );
AOI21X1 AOI21X1_928 ( .A(reg_pc_5_), .B(decoded_imm_5_), .C(_2516_), .Y(_2517_) );
OAI21X1 OAI21X1_3331 ( .A(_2485_), .B(_2515_), .C(_2517_), .Y(_2518_) );
NAND2X1 NAND2X1_1015 ( .A(_4658_), .B(_8005_), .Y(_2519_) );
NOR2X1 NOR2X1_1250 ( .A(_4658_), .B(_8005_), .Y(_2520_) );
INVX1 INVX1_1194 ( .A(_2520_), .Y(_2521_) );
NAND2X1 NAND2X1_1016 ( .A(_2519_), .B(_2521_), .Y(_2522_) );
INVX1 INVX1_1195 ( .A(_2522_), .Y(_2523_) );
AND2X2 AND2X2_202 ( .A(_2518_), .B(_2523_), .Y(_2524_) );
OAI21X1 OAI21X1_3332 ( .A(_2518_), .B(_2523_), .C(cpu_state_3_bF_buf3_), .Y(_2525_) );
NAND2X1 NAND2X1_1017 ( .A(mem_rdata[30]), .B(_2414_), .Y(_2526_) );
OAI21X1 OAI21X1_3333 ( .A(_2467_), .B(_4617_), .C(_2526_), .Y(_2527_) );
NAND2X1 NAND2X1_1018 ( .A(_1816_), .B(_2527_), .Y(_2528_) );
AOI22X1 AOI22X1_139 ( .A(mem_rdata[22]), .B(_1809_), .C(_10730__0_), .D(mem_rdata[6]), .Y(_2529_) );
AOI21X1 AOI21X1_929 ( .A(_2528_), .B(_2529_), .C(_4448_), .Y(_2530_) );
AND2X2 AND2X2_203 ( .A(_2421_), .B(count_instr_38_), .Y(_2531_) );
AOI22X1 AOI22X1_140 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_6_), .C(instr_rdcycleh_bF_buf1), .D(count_cycle_38_), .Y(_2532_) );
OAI21X1 OAI21X1_3334 ( .A(_4529_), .B(_1238_), .C(_2532_), .Y(_2533_) );
OAI21X1 OAI21X1_3335 ( .A(_2531_), .B(_2533_), .C(cpu_state_2_bF_buf5_), .Y(_2534_) );
OAI21X1 OAI21X1_3336 ( .A(_4575__bF_buf1), .B(_5174_), .C(_2534_), .Y(_2535_) );
NOR2X1 NOR2X1_1251 ( .A(_2530_), .B(_2535_), .Y(_2536_) );
OAI21X1 OAI21X1_3337 ( .A(_2524_), .B(_2525_), .C(_2536_), .Y(_83__6_) );
XNOR2X1 XNOR2X1_54 ( .A(reg_pc_7_), .B(decoded_imm_7_), .Y(_2537_) );
NOR2X1 NOR2X1_1252 ( .A(_2520_), .B(_2524_), .Y(_2538_) );
XOR2X1 XOR2X1_9 ( .A(_2538_), .B(_2537_), .Y(_2539_) );
NAND2X1 NAND2X1_1019 ( .A(mem_rdata[31]), .B(_2414_), .Y(_2540_) );
OAI21X1 OAI21X1_3338 ( .A(_2467_), .B(_1535_), .C(_2540_), .Y(_2541_) );
OAI21X1 OAI21X1_3339 ( .A(_1798_), .B(_2465_), .C(mem_rdata[7]), .Y(_2542_) );
OAI21X1 OAI21X1_3340 ( .A(_1810_), .B(_1513_), .C(_2542_), .Y(_2543_) );
AOI21X1 AOI21X1_930 ( .A(_1816_), .B(_2541_), .C(_2543_), .Y(_2544_) );
INVX1 INVX1_1196 ( .A(count_cycle_39_), .Y(_2545_) );
NOR2X1 NOR2X1_1253 ( .A(_1735_), .B(_2545_), .Y(_2546_) );
AOI22X1 AOI22X1_141 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_7_), .C(instr_rdinstr_bF_buf3), .D(count_instr_7_), .Y(_2547_) );
OAI21X1 OAI21X1_3341 ( .A(_4531__bF_buf2), .B(_1380_), .C(_2547_), .Y(_2548_) );
OAI21X1 OAI21X1_3342 ( .A(_2548_), .B(_2546_), .C(cpu_state_2_bF_buf4_), .Y(_2549_) );
OAI21X1 OAI21X1_3343 ( .A(_2544_), .B(_4448_), .C(_2549_), .Y(_2550_) );
AOI21X1 AOI21X1_931 ( .A(cpu_state_3_bF_buf2_), .B(_2539_), .C(_2550_), .Y(_2551_) );
OAI21X1 OAI21X1_3344 ( .A(_4575__bF_buf0), .B(_5173_), .C(_2551_), .Y(_83__7_) );
NOR2X1 NOR2X1_1254 ( .A(_2537_), .B(_2522_), .Y(_2552_) );
INVX1 INVX1_1197 ( .A(_2552_), .Y(_2553_) );
NOR2X1 NOR2X1_1255 ( .A(_2537_), .B(_2521_), .Y(_2554_) );
AOI21X1 AOI21X1_932 ( .A(reg_pc_7_), .B(decoded_imm_7_), .C(_2554_), .Y(_2555_) );
OAI21X1 OAI21X1_3345 ( .A(_2553_), .B(_2517_), .C(_2555_), .Y(_2556_) );
INVX1 INVX1_1198 ( .A(_2556_), .Y(_2557_) );
NAND2X1 NAND2X1_1020 ( .A(_2514_), .B(_2552_), .Y(_2558_) );
OAI21X1 OAI21X1_3346 ( .A(_2485_), .B(_2558_), .C(_2557_), .Y(_2559_) );
NAND2X1 NAND2X1_1021 ( .A(_4679_), .B(_8230_), .Y(_2560_) );
NOR2X1 NOR2X1_1256 ( .A(_4679_), .B(_8230_), .Y(_2561_) );
INVX1 INVX1_1199 ( .A(_2561_), .Y(_2562_) );
AND2X2 AND2X2_204 ( .A(_2562_), .B(_2560_), .Y(_2563_) );
NOR2X1 NOR2X1_1257 ( .A(_2563_), .B(_2559_), .Y(_2564_) );
NAND2X1 NAND2X1_1022 ( .A(_2563_), .B(_2559_), .Y(_2565_) );
NAND2X1 NAND2X1_1023 ( .A(cpu_state_3_bF_buf1_), .B(_2565_), .Y(_2566_) );
INVX1 INVX1_1200 ( .A(latched_is_lu), .Y(_2567_) );
INVX1 INVX1_1201 ( .A(latched_is_lh), .Y(_2568_) );
NAND2X1 NAND2X1_1024 ( .A(_2567_), .B(_2568_), .Y(_2569_) );
OAI22X1 OAI22X1_276 ( .A(_1529_), .B(_1808_), .C(_1799_), .D(_1693_), .Y(_2570_) );
NOR2X1 NOR2X1_1258 ( .A(_2569_), .B(_2544_), .Y(_2571_) );
AOI21X1 AOI21X1_933 ( .A(_2569_), .B(_2570_), .C(_2571_), .Y(_2572_) );
NOR2X1 NOR2X1_1259 ( .A(_1393_), .B(_4531__bF_buf1), .Y(_2573_) );
NAND2X1 NAND2X1_1025 ( .A(instr_rdinstr_bF_buf2), .B(count_instr_8_), .Y(_2574_) );
NAND2X1 NAND2X1_1026 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_8_), .Y(_2575_) );
NAND2X1 NAND2X1_1027 ( .A(instr_rdcycleh_bF_buf0), .B(count_cycle_40_), .Y(_2576_) );
NAND3X1 NAND3X1_98 ( .A(_2574_), .B(_2575_), .C(_2576_), .Y(_2577_) );
OAI21X1 OAI21X1_3347 ( .A(_2573_), .B(_2577_), .C(cpu_state_2_bF_buf3_), .Y(_2578_) );
OAI21X1 OAI21X1_3348 ( .A(_2572_), .B(_4448_), .C(_2578_), .Y(_2579_) );
AOI21X1 AOI21X1_934 ( .A(cpu_state_4_), .B(_10734__8_), .C(_2579_), .Y(_2580_) );
OAI21X1 OAI21X1_3349 ( .A(_2566_), .B(_2564_), .C(_2580_), .Y(_83__8_) );
OAI22X1 OAI22X1_277 ( .A(_1516_), .B(_1808_), .C(_1799_), .D(_1696_), .Y(_2581_) );
AOI21X1 AOI21X1_935 ( .A(_2569_), .B(_2581_), .C(_2571_), .Y(_2582_) );
NOR2X1 NOR2X1_1260 ( .A(reg_pc_9_), .B(decoded_imm_9_), .Y(_2583_) );
NOR2X1 NOR2X1_1261 ( .A(_8237_), .B(_8225_), .Y(_2584_) );
OR2X2 OR2X2_42 ( .A(_2584_), .B(_2583_), .Y(_2585_) );
INVX1 INVX1_1202 ( .A(_2585_), .Y(_2586_) );
NOR2X1 NOR2X1_1262 ( .A(_2561_), .B(_2586_), .Y(_2587_) );
AOI21X1 AOI21X1_936 ( .A(_2562_), .B(_2565_), .C(_2585_), .Y(_2588_) );
AOI21X1 AOI21X1_937 ( .A(_2565_), .B(_2587_), .C(_2588_), .Y(_2589_) );
NOR2X1 NOR2X1_1263 ( .A(_1388_), .B(_4531__bF_buf0), .Y(_2590_) );
INVX1 INVX1_1203 ( .A(count_cycle_41_), .Y(_2591_) );
AOI22X1 AOI22X1_142 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_9_), .C(instr_rdinstr_bF_buf1), .D(count_instr_9_), .Y(_2592_) );
OAI21X1 OAI21X1_3350 ( .A(_1735_), .B(_2591_), .C(_2592_), .Y(_2593_) );
OAI21X1 OAI21X1_3351 ( .A(_2590_), .B(_2593_), .C(cpu_state_2_bF_buf2_), .Y(_2594_) );
OAI21X1 OAI21X1_3352 ( .A(_4575__bF_buf4), .B(_5107_), .C(_2594_), .Y(_2595_) );
AOI21X1 AOI21X1_938 ( .A(cpu_state_3_bF_buf0_), .B(_2589_), .C(_2595_), .Y(_2596_) );
OAI21X1 OAI21X1_3353 ( .A(_4448_), .B(_2582_), .C(_2596_), .Y(_83__9_) );
INVX1 INVX1_1204 ( .A(_2559_), .Y(_2597_) );
NAND2X1 NAND2X1_1028 ( .A(_2563_), .B(_2586_), .Y(_2598_) );
NOR2X1 NOR2X1_1264 ( .A(_2562_), .B(_2585_), .Y(_2599_) );
NOR2X1 NOR2X1_1265 ( .A(_2584_), .B(_2599_), .Y(_2600_) );
OAI21X1 OAI21X1_3354 ( .A(_2597_), .B(_2598_), .C(_2600_), .Y(_2601_) );
NOR2X1 NOR2X1_1266 ( .A(reg_pc_10_), .B(decoded_imm_10_), .Y(_2602_) );
NAND2X1 NAND2X1_1029 ( .A(reg_pc_10_), .B(decoded_imm_10_), .Y(_2603_) );
INVX1 INVX1_1205 ( .A(_2603_), .Y(_2604_) );
NOR2X1 NOR2X1_1267 ( .A(_2602_), .B(_2604_), .Y(_2605_) );
NOR2X1 NOR2X1_1268 ( .A(_2605_), .B(_2601_), .Y(_2606_) );
NOR2X1 NOR2X1_1269 ( .A(_2598_), .B(_2597_), .Y(_2607_) );
INVX1 INVX1_1206 ( .A(_2600_), .Y(_2608_) );
OAI21X1 OAI21X1_3355 ( .A(_2607_), .B(_2608_), .C(_2605_), .Y(_2609_) );
NAND2X1 NAND2X1_1030 ( .A(cpu_state_3_bF_buf4_), .B(_2609_), .Y(_2610_) );
OAI22X1 OAI22X1_278 ( .A(_1504_), .B(_1808_), .C(_1799_), .D(_1699_), .Y(_2611_) );
AOI21X1 AOI21X1_939 ( .A(_2569_), .B(_2611_), .C(_2571_), .Y(_2612_) );
NOR2X1 NOR2X1_1270 ( .A(_1397_), .B(_4531__bF_buf4), .Y(_2613_) );
NAND2X1 NAND2X1_1031 ( .A(instr_rdinstr_bF_buf0), .B(count_instr_10_), .Y(_2614_) );
NAND2X1 NAND2X1_1032 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_10_), .Y(_2615_) );
NAND2X1 NAND2X1_1033 ( .A(instr_rdcycleh_bF_buf3), .B(count_cycle_42_), .Y(_2616_) );
NAND3X1 NAND3X1_99 ( .A(_2614_), .B(_2615_), .C(_2616_), .Y(_2617_) );
OAI21X1 OAI21X1_3356 ( .A(_2613_), .B(_2617_), .C(cpu_state_2_bF_buf1_), .Y(_2618_) );
OAI21X1 OAI21X1_3357 ( .A(_2612_), .B(_4448_), .C(_2618_), .Y(_2619_) );
AOI21X1 AOI21X1_940 ( .A(cpu_state_4_), .B(_10734__10_), .C(_2619_), .Y(_2620_) );
OAI21X1 OAI21X1_3358 ( .A(_2610_), .B(_2606_), .C(_2620_), .Y(_83__10_) );
NAND2X1 NAND2X1_1034 ( .A(_2603_), .B(_2609_), .Y(_2621_) );
NOR2X1 NOR2X1_1271 ( .A(reg_pc_11_), .B(decoded_imm_11_), .Y(_2622_) );
NAND2X1 NAND2X1_1035 ( .A(reg_pc_11_), .B(decoded_imm_11_), .Y(_2623_) );
INVX1 INVX1_1207 ( .A(_2623_), .Y(_2624_) );
NOR2X1 NOR2X1_1272 ( .A(_2622_), .B(_2624_), .Y(_2625_) );
XNOR2X1 XNOR2X1_55 ( .A(_2621_), .B(_2625_), .Y(_2626_) );
OAI22X1 OAI22X1_279 ( .A(_1501_), .B(_1808_), .C(_1799_), .D(_1702_), .Y(_2627_) );
AOI21X1 AOI21X1_941 ( .A(_2569_), .B(_2627_), .C(_2571_), .Y(_2628_) );
NOR2X1 NOR2X1_1273 ( .A(_1402_), .B(_4531__bF_buf3), .Y(_2629_) );
NAND2X1 NAND2X1_1036 ( .A(instr_rdinstr_bF_buf4), .B(count_instr_11_), .Y(_2630_) );
NAND2X1 NAND2X1_1037 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_11_), .Y(_2631_) );
NAND2X1 NAND2X1_1038 ( .A(instr_rdcycleh_bF_buf2), .B(count_cycle_43_), .Y(_2632_) );
NAND3X1 NAND3X1_100 ( .A(_2630_), .B(_2631_), .C(_2632_), .Y(_2633_) );
OAI21X1 OAI21X1_3359 ( .A(_2629_), .B(_2633_), .C(cpu_state_2_bF_buf0_), .Y(_2634_) );
OAI21X1 OAI21X1_3360 ( .A(_2628_), .B(_4448_), .C(_2634_), .Y(_2635_) );
AOI21X1 AOI21X1_942 ( .A(cpu_state_4_), .B(_10734__11_), .C(_2635_), .Y(_2636_) );
OAI21X1 OAI21X1_3361 ( .A(_2626_), .B(_4555_), .C(_2636_), .Y(_83__11_) );
NAND2X1 NAND2X1_1039 ( .A(_2605_), .B(_2625_), .Y(_2637_) );
NOR2X1 NOR2X1_1274 ( .A(_2637_), .B(_2598_), .Y(_2638_) );
INVX1 INVX1_1208 ( .A(_2638_), .Y(_2639_) );
INVX1 INVX1_1209 ( .A(_2637_), .Y(_2640_) );
OAI21X1 OAI21X1_3362 ( .A(_2622_), .B(_2603_), .C(_2623_), .Y(_2641_) );
AOI21X1 AOI21X1_943 ( .A(_2640_), .B(_2608_), .C(_2641_), .Y(_2642_) );
OAI21X1 OAI21X1_3363 ( .A(_2597_), .B(_2639_), .C(_2642_), .Y(_2643_) );
NAND2X1 NAND2X1_1040 ( .A(_4719_), .B(_8465_), .Y(_2644_) );
NOR2X1 NOR2X1_1275 ( .A(_4719_), .B(_8465_), .Y(_2645_) );
INVX1 INVX1_1210 ( .A(_2645_), .Y(_2646_) );
AND2X2 AND2X2_205 ( .A(_2646_), .B(_2644_), .Y(_2647_) );
NOR2X1 NOR2X1_1276 ( .A(_2647_), .B(_2643_), .Y(_2648_) );
INVX1 INVX1_1211 ( .A(_2643_), .Y(_2649_) );
INVX1 INVX1_1212 ( .A(_2647_), .Y(_2650_) );
OAI21X1 OAI21X1_3364 ( .A(_2649_), .B(_2650_), .C(cpu_state_3_bF_buf3_), .Y(_2651_) );
OAI22X1 OAI22X1_280 ( .A(_1519_), .B(_1808_), .C(_1799_), .D(_4613_), .Y(_2652_) );
AOI21X1 AOI21X1_944 ( .A(_2569_), .B(_2652_), .C(_2571_), .Y(_2653_) );
NOR2X1 NOR2X1_1277 ( .A(_1407_), .B(_4531__bF_buf2), .Y(_2654_) );
NAND2X1 NAND2X1_1041 ( .A(instr_rdinstr_bF_buf3), .B(count_instr_12_), .Y(_2655_) );
NAND2X1 NAND2X1_1042 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_12_), .Y(_2656_) );
NAND2X1 NAND2X1_1043 ( .A(instr_rdcycleh_bF_buf1), .B(count_cycle_44_), .Y(_2657_) );
NAND3X1 NAND3X1_101 ( .A(_2655_), .B(_2656_), .C(_2657_), .Y(_2658_) );
OAI21X1 OAI21X1_3365 ( .A(_2654_), .B(_2658_), .C(cpu_state_2_bF_buf5_), .Y(_2659_) );
OAI21X1 OAI21X1_3366 ( .A(_2653_), .B(_4448_), .C(_2659_), .Y(_2660_) );
AOI21X1 AOI21X1_945 ( .A(cpu_state_4_), .B(_10734__12_), .C(_2660_), .Y(_2661_) );
OAI21X1 OAI21X1_3367 ( .A(_2651_), .B(_2648_), .C(_2661_), .Y(_83__12_) );
OAI22X1 OAI22X1_281 ( .A(_1522_), .B(_1808_), .C(_1799_), .D(_4615_), .Y(_2662_) );
AOI21X1 AOI21X1_946 ( .A(_2569_), .B(_2662_), .C(_2571_), .Y(_2663_) );
NOR2X1 NOR2X1_1278 ( .A(reg_pc_13_), .B(decoded_imm_13_), .Y(_2664_) );
NOR2X1 NOR2X1_1279 ( .A(_4768_), .B(_8543_), .Y(_2665_) );
NOR2X1 NOR2X1_1280 ( .A(_2664_), .B(_2665_), .Y(_2666_) );
OAI21X1 OAI21X1_3368 ( .A(_2649_), .B(_2650_), .C(_2646_), .Y(_2667_) );
XOR2X1 XOR2X1_10 ( .A(_2667_), .B(_2666_), .Y(_2668_) );
NOR2X1 NOR2X1_1281 ( .A(_1412_), .B(_4531__bF_buf1), .Y(_2669_) );
AOI22X1 AOI22X1_143 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_13_), .C(instr_rdcycleh_bF_buf0), .D(count_cycle_45_), .Y(_2670_) );
OAI21X1 OAI21X1_3369 ( .A(_4529_), .B(_1270_), .C(_2670_), .Y(_2671_) );
OAI21X1 OAI21X1_3370 ( .A(_2669_), .B(_2671_), .C(cpu_state_2_bF_buf4_), .Y(_2672_) );
OAI21X1 OAI21X1_3371 ( .A(_4575__bF_buf3), .B(_5196_), .C(_2672_), .Y(_2673_) );
AOI21X1 AOI21X1_947 ( .A(cpu_state_3_bF_buf2_), .B(_2668_), .C(_2673_), .Y(_2674_) );
OAI21X1 OAI21X1_3372 ( .A(_4448_), .B(_2663_), .C(_2674_), .Y(_83__13_) );
NAND2X1 NAND2X1_1044 ( .A(_2666_), .B(_2647_), .Y(_2675_) );
NOR2X1 NOR2X1_1282 ( .A(_2675_), .B(_2649_), .Y(_2676_) );
INVX1 INVX1_1213 ( .A(_2665_), .Y(_2677_) );
OAI21X1 OAI21X1_3373 ( .A(_2646_), .B(_2664_), .C(_2677_), .Y(_2678_) );
NAND2X1 NAND2X1_1045 ( .A(_4736_), .B(_8623_), .Y(_2679_) );
NOR2X1 NOR2X1_1283 ( .A(_4736_), .B(_8623_), .Y(_2680_) );
INVX1 INVX1_1214 ( .A(_2680_), .Y(_2681_) );
AND2X2 AND2X2_206 ( .A(_2681_), .B(_2679_), .Y(_2682_) );
OAI21X1 OAI21X1_3374 ( .A(_2676_), .B(_2678_), .C(_2682_), .Y(_2683_) );
NOR2X1 NOR2X1_1284 ( .A(_2678_), .B(_2676_), .Y(_2684_) );
INVX1 INVX1_1215 ( .A(_2682_), .Y(_2685_) );
NAND2X1 NAND2X1_1046 ( .A(_2685_), .B(_2684_), .Y(_2686_) );
NAND2X1 NAND2X1_1047 ( .A(_2683_), .B(_2686_), .Y(_2687_) );
OAI22X1 OAI22X1_282 ( .A(_1498_), .B(_1808_), .C(_1799_), .D(_4617_), .Y(_2688_) );
AOI21X1 AOI21X1_948 ( .A(_2569_), .B(_2688_), .C(_2571_), .Y(_2689_) );
NOR2X1 NOR2X1_1285 ( .A(_1425_), .B(_4531__bF_buf0), .Y(_2690_) );
INVX1 INVX1_1216 ( .A(count_cycle_46_), .Y(_2691_) );
AOI22X1 AOI22X1_144 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_14_), .C(instr_rdinstr_bF_buf2), .D(count_instr_14_), .Y(_2692_) );
OAI21X1 OAI21X1_3375 ( .A(_1735_), .B(_2691_), .C(_2692_), .Y(_2693_) );
OAI21X1 OAI21X1_3376 ( .A(_2690_), .B(_2693_), .C(cpu_state_2_bF_buf3_), .Y(_2694_) );
OAI21X1 OAI21X1_3377 ( .A(_2689_), .B(_4448_), .C(_2694_), .Y(_2695_) );
AOI21X1 AOI21X1_949 ( .A(cpu_state_4_), .B(_10734__14_), .C(_2695_), .Y(_2696_) );
OAI21X1 OAI21X1_3378 ( .A(_2687_), .B(_4555_), .C(_2696_), .Y(_83__14_) );
OAI21X1 OAI21X1_3379 ( .A(_4736_), .B(_8623_), .C(_2683_), .Y(_2697_) );
NOR2X1 NOR2X1_1286 ( .A(reg_pc_15_), .B(decoded_imm_15_), .Y(_2698_) );
NAND2X1 NAND2X1_1048 ( .A(reg_pc_15_), .B(decoded_imm_15_), .Y(_2699_) );
INVX1 INVX1_1217 ( .A(_2699_), .Y(_2700_) );
NOR2X1 NOR2X1_1287 ( .A(_2698_), .B(_2700_), .Y(_2701_) );
AND2X2 AND2X2_207 ( .A(_2697_), .B(_2701_), .Y(_2702_) );
OAI21X1 OAI21X1_3380 ( .A(_2697_), .B(_2701_), .C(cpu_state_3_bF_buf1_), .Y(_2703_) );
OAI22X1 OAI22X1_283 ( .A(_1525_), .B(_1808_), .C(_1799_), .D(_1535_), .Y(_2704_) );
AOI21X1 AOI21X1_950 ( .A(_2569_), .B(_2704_), .C(_2571_), .Y(_2705_) );
INVX1 INVX1_1218 ( .A(count_cycle_47_), .Y(_2706_) );
NOR2X1 NOR2X1_1288 ( .A(_1735_), .B(_2706_), .Y(_2707_) );
AOI22X1 AOI22X1_145 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_15_), .C(instr_rdinstr_bF_buf1), .D(count_instr_15_), .Y(_2708_) );
OAI21X1 OAI21X1_3381 ( .A(_4531__bF_buf4), .B(_1422_), .C(_2708_), .Y(_2709_) );
OAI21X1 OAI21X1_3382 ( .A(_2709_), .B(_2707_), .C(cpu_state_2_bF_buf2_), .Y(_2710_) );
OAI21X1 OAI21X1_3383 ( .A(_2705_), .B(_4448_), .C(_2710_), .Y(_2711_) );
AOI21X1 AOI21X1_951 ( .A(cpu_state_4_), .B(_10734__15_), .C(_2711_), .Y(_2712_) );
OAI21X1 OAI21X1_3384 ( .A(_2702_), .B(_2703_), .C(_2712_), .Y(_83__15_) );
NAND2X1 NAND2X1_1049 ( .A(_2701_), .B(_2682_), .Y(_2713_) );
NOR2X1 NOR2X1_1289 ( .A(_2675_), .B(_2713_), .Y(_2714_) );
INVX1 INVX1_1219 ( .A(_2714_), .Y(_2715_) );
NAND3X1 NAND3X1_102 ( .A(_2701_), .B(_2678_), .C(_2682_), .Y(_2716_) );
AOI21X1 AOI21X1_952 ( .A(_2680_), .B(_2701_), .C(_2700_), .Y(_2717_) );
AND2X2 AND2X2_208 ( .A(_2716_), .B(_2717_), .Y(_2718_) );
OAI21X1 OAI21X1_3385 ( .A(_2642_), .B(_2715_), .C(_2718_), .Y(_2719_) );
NAND2X1 NAND2X1_1050 ( .A(_2714_), .B(_2638_), .Y(_2720_) );
NOR2X1 NOR2X1_1290 ( .A(_2720_), .B(_2597_), .Y(_2721_) );
OR2X2 OR2X2_43 ( .A(_2721_), .B(_2719_), .Y(_2722_) );
NAND2X1 NAND2X1_1051 ( .A(_4774_), .B(_8782_), .Y(_2723_) );
NOR2X1 NOR2X1_1291 ( .A(_4774_), .B(_8782_), .Y(_2724_) );
INVX1 INVX1_1220 ( .A(_2724_), .Y(_2725_) );
AND2X2 AND2X2_209 ( .A(_2725_), .B(_2723_), .Y(_2726_) );
NOR2X1 NOR2X1_1292 ( .A(_2726_), .B(_2722_), .Y(_2727_) );
NOR2X1 NOR2X1_1293 ( .A(_2719_), .B(_2721_), .Y(_2728_) );
INVX1 INVX1_1221 ( .A(_2726_), .Y(_2729_) );
OAI21X1 OAI21X1_3386 ( .A(_2728_), .B(_2729_), .C(cpu_state_3_bF_buf0_), .Y(_2730_) );
NOR2X1 NOR2X1_1294 ( .A(_4425_), .B(_2567_), .Y(_2731_) );
AND2X2 AND2X2_210 ( .A(_2704_), .B(latched_is_lh), .Y(_2732_) );
AOI21X1 AOI21X1_953 ( .A(mem_rdata[16]), .B(_2731_), .C(_2732_), .Y(_2733_) );
OAI21X1 OAI21X1_3387 ( .A(_2544_), .B(_2569_), .C(_2733_), .Y(_2734_) );
NOR2X1 NOR2X1_1295 ( .A(_1432_), .B(_4531__bF_buf3), .Y(_2735_) );
AOI22X1 AOI22X1_146 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_16_), .C(instr_rdcycleh_bF_buf3), .D(count_cycle_48_), .Y(_2736_) );
OAI21X1 OAI21X1_3388 ( .A(_4529_), .B(_1278_), .C(_2736_), .Y(_2737_) );
OAI21X1 OAI21X1_3389 ( .A(_2735_), .B(_2737_), .C(cpu_state_2_bF_buf1_), .Y(_2738_) );
OAI21X1 OAI21X1_3390 ( .A(_4575__bF_buf2), .B(_5051_), .C(_2738_), .Y(_2739_) );
AOI21X1 AOI21X1_954 ( .A(_4447__bF_buf0), .B(_2734_), .C(_2739_), .Y(_2740_) );
OAI21X1 OAI21X1_3391 ( .A(_2727_), .B(_2730_), .C(_2740_), .Y(_83__16_) );
NOR2X1 NOR2X1_1296 ( .A(reg_pc_17_), .B(decoded_imm_17_), .Y(_2741_) );
NOR2X1 NOR2X1_1297 ( .A(_4775_), .B(_8868_), .Y(_2742_) );
NOR2X1 NOR2X1_1298 ( .A(_2741_), .B(_2742_), .Y(_2743_) );
INVX1 INVX1_1222 ( .A(_2743_), .Y(_2744_) );
NOR2X1 NOR2X1_1299 ( .A(_2744_), .B(_2729_), .Y(_2745_) );
OAI21X1 OAI21X1_3392 ( .A(_2721_), .B(_2719_), .C(_2745_), .Y(_2746_) );
INVX1 INVX1_1223 ( .A(_2746_), .Y(_2747_) );
OAI21X1 OAI21X1_3393 ( .A(_2721_), .B(_2719_), .C(_2726_), .Y(_2748_) );
OAI21X1 OAI21X1_3394 ( .A(_4774_), .B(_8782_), .C(_2748_), .Y(_2749_) );
NOR2X1 NOR2X1_1300 ( .A(_2725_), .B(_2744_), .Y(_2750_) );
NOR2X1 NOR2X1_1301 ( .A(_4555_), .B(_2750_), .Y(_2751_) );
OAI21X1 OAI21X1_3395 ( .A(_2749_), .B(_2743_), .C(_2751_), .Y(_2752_) );
NAND2X1 NAND2X1_1052 ( .A(mem_wordsize_0_bF_buf0_), .B(latched_is_lu), .Y(_2753_) );
NOR2X1 NOR2X1_1302 ( .A(_2732_), .B(_2571_), .Y(_2754_) );
OAI21X1 OAI21X1_3396 ( .A(_1541_), .B(_2753_), .C(_2754_), .Y(_2755_) );
INVX1 INVX1_1224 ( .A(count_cycle_49_), .Y(_2756_) );
NOR2X1 NOR2X1_1303 ( .A(_1735_), .B(_2756_), .Y(_2757_) );
AOI22X1 AOI22X1_147 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_17_), .C(instr_rdinstr_bF_buf0), .D(count_instr_17_), .Y(_2758_) );
OAI21X1 OAI21X1_3397 ( .A(_4531__bF_buf2), .B(_1433_), .C(_2758_), .Y(_2759_) );
OAI21X1 OAI21X1_3398 ( .A(_2759_), .B(_2757_), .C(cpu_state_2_bF_buf0_), .Y(_2760_) );
OAI21X1 OAI21X1_3399 ( .A(_4575__bF_buf1), .B(_5057_), .C(_2760_), .Y(_2761_) );
AOI21X1 AOI21X1_955 ( .A(_4447__bF_buf3), .B(_2755_), .C(_2761_), .Y(_2762_) );
OAI21X1 OAI21X1_3400 ( .A(_2752_), .B(_2747_), .C(_2762_), .Y(_83__17_) );
NOR2X1 NOR2X1_1304 ( .A(_2742_), .B(_2750_), .Y(_2763_) );
OAI21X1 OAI21X1_3401 ( .A(_2748_), .B(_2744_), .C(_2763_), .Y(_2764_) );
NOR2X1 NOR2X1_1305 ( .A(reg_pc_18_), .B(decoded_imm_18_), .Y(_2765_) );
NOR2X1 NOR2X1_1306 ( .A(_4779_), .B(_8947_), .Y(_2766_) );
NOR2X1 NOR2X1_1307 ( .A(_2765_), .B(_2766_), .Y(_2767_) );
XNOR2X1 XNOR2X1_56 ( .A(_2764_), .B(_2767_), .Y(_2768_) );
OAI21X1 OAI21X1_3402 ( .A(_1544_), .B(_2753_), .C(_2754_), .Y(_2769_) );
NOR2X1 NOR2X1_1308 ( .A(_1437_), .B(_4531__bF_buf1), .Y(_2770_) );
NAND2X1 NAND2X1_1053 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_18_), .Y(_2771_) );
NAND2X1 NAND2X1_1054 ( .A(instr_rdinstr_bF_buf4), .B(count_instr_18_), .Y(_2772_) );
NAND2X1 NAND2X1_1055 ( .A(instr_rdcycleh_bF_buf2), .B(count_cycle_50_), .Y(_2773_) );
NAND3X1 NAND3X1_103 ( .A(_2771_), .B(_2772_), .C(_2773_), .Y(_2774_) );
OAI21X1 OAI21X1_3403 ( .A(_2770_), .B(_2774_), .C(cpu_state_2_bF_buf5_), .Y(_2775_) );
OAI21X1 OAI21X1_3404 ( .A(_4575__bF_buf0), .B(_5045_), .C(_2775_), .Y(_2776_) );
AOI21X1 AOI21X1_956 ( .A(_4447__bF_buf2), .B(_2769_), .C(_2776_), .Y(_2777_) );
OAI21X1 OAI21X1_3405 ( .A(_2768_), .B(_4555_), .C(_2777_), .Y(_83__18_) );
AOI21X1 AOI21X1_957 ( .A(_2767_), .B(_2764_), .C(_2766_), .Y(_2778_) );
NOR2X1 NOR2X1_1309 ( .A(reg_pc_19_), .B(decoded_imm_19_), .Y(_2779_) );
NOR2X1 NOR2X1_1310 ( .A(_4790_), .B(_1647_), .Y(_2780_) );
NOR2X1 NOR2X1_1311 ( .A(_2779_), .B(_2780_), .Y(_2781_) );
INVX1 INVX1_1225 ( .A(_2781_), .Y(_2782_) );
AND2X2 AND2X2_211 ( .A(_2778_), .B(_2782_), .Y(_2783_) );
OAI21X1 OAI21X1_3406 ( .A(_2778_), .B(_2782_), .C(cpu_state_3_bF_buf4_), .Y(_2784_) );
OAI21X1 OAI21X1_3407 ( .A(_1495_), .B(_2753_), .C(_2754_), .Y(_2785_) );
INVX1 INVX1_1226 ( .A(count_cycle_51_), .Y(_2786_) );
NOR2X1 NOR2X1_1312 ( .A(_1735_), .B(_2786_), .Y(_2787_) );
AOI22X1 AOI22X1_148 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_19_), .C(instr_rdinstr_bF_buf3), .D(count_instr_19_), .Y(_2788_) );
OAI21X1 OAI21X1_3408 ( .A(_4531__bF_buf0), .B(_1445_), .C(_2788_), .Y(_2789_) );
OAI21X1 OAI21X1_3409 ( .A(_2789_), .B(_2787_), .C(cpu_state_2_bF_buf4_), .Y(_2790_) );
OAI21X1 OAI21X1_3410 ( .A(_4575__bF_buf4), .B(_5040_), .C(_2790_), .Y(_2791_) );
AOI21X1 AOI21X1_958 ( .A(_4447__bF_buf1), .B(_2785_), .C(_2791_), .Y(_2792_) );
OAI21X1 OAI21X1_3411 ( .A(_2783_), .B(_2784_), .C(_2792_), .Y(_83__19_) );
NAND2X1 NAND2X1_1056 ( .A(_2781_), .B(_2767_), .Y(_2793_) );
INVX1 INVX1_1227 ( .A(_2793_), .Y(_2794_) );
NAND2X1 NAND2X1_1057 ( .A(_2794_), .B(_2745_), .Y(_2795_) );
INVX1 INVX1_1228 ( .A(_2795_), .Y(_2796_) );
AOI21X1 AOI21X1_959 ( .A(_2766_), .B(_2781_), .C(_2780_), .Y(_2797_) );
OAI21X1 OAI21X1_3412 ( .A(_2763_), .B(_2793_), .C(_2797_), .Y(_2798_) );
AOI21X1 AOI21X1_960 ( .A(_2796_), .B(_2722_), .C(_2798_), .Y(_2799_) );
NOR2X1 NOR2X1_1313 ( .A(reg_pc_20_), .B(decoded_imm_20_), .Y(_2800_) );
NOR2X1 NOR2X1_1314 ( .A(_4803_), .B(_9107_), .Y(_2801_) );
NOR2X1 NOR2X1_1315 ( .A(_2800_), .B(_2801_), .Y(_2802_) );
INVX1 INVX1_1229 ( .A(_2802_), .Y(_2803_) );
AND2X2 AND2X2_212 ( .A(_2799_), .B(_2803_), .Y(_2804_) );
OAI21X1 OAI21X1_3413 ( .A(_2799_), .B(_2803_), .C(cpu_state_3_bF_buf3_), .Y(_2805_) );
OAI21X1 OAI21X1_3414 ( .A(_1532_), .B(_2753_), .C(_2754_), .Y(_2806_) );
NOR2X1 NOR2X1_1316 ( .A(_1449_), .B(_4531__bF_buf4), .Y(_2807_) );
AOI22X1 AOI22X1_149 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_20_), .C(instr_rdcycleh_bF_buf1), .D(count_cycle_52_), .Y(_2808_) );
OAI21X1 OAI21X1_3415 ( .A(_4529_), .B(_1297_), .C(_2808_), .Y(_2809_) );
OAI21X1 OAI21X1_3416 ( .A(_2807_), .B(_2809_), .C(cpu_state_2_bF_buf3_), .Y(_2810_) );
OAI21X1 OAI21X1_3417 ( .A(_4575__bF_buf3), .B(_5218_), .C(_2810_), .Y(_2811_) );
AOI21X1 AOI21X1_961 ( .A(_4447__bF_buf0), .B(_2806_), .C(_2811_), .Y(_2812_) );
OAI21X1 OAI21X1_3418 ( .A(_2804_), .B(_2805_), .C(_2812_), .Y(_83__20_) );
NOR2X1 NOR2X1_1317 ( .A(reg_pc_21_), .B(decoded_imm_21_), .Y(_2813_) );
NOR2X1 NOR2X1_1318 ( .A(_4812_), .B(_1654_), .Y(_2814_) );
NOR2X1 NOR2X1_1319 ( .A(_2813_), .B(_2814_), .Y(_2815_) );
INVX1 INVX1_1230 ( .A(_2815_), .Y(_2816_) );
INVX1 INVX1_1231 ( .A(_2799_), .Y(_2817_) );
AOI21X1 AOI21X1_962 ( .A(_2802_), .B(_2817_), .C(_2801_), .Y(_2818_) );
AND2X2 AND2X2_213 ( .A(_2818_), .B(_2816_), .Y(_2819_) );
OAI21X1 OAI21X1_3419 ( .A(_2818_), .B(_2816_), .C(cpu_state_3_bF_buf2_), .Y(_2820_) );
OAI21X1 OAI21X1_3420 ( .A(_2500_), .B(_2753_), .C(_2754_), .Y(_2821_) );
NOR2X1 NOR2X1_1320 ( .A(_1451_), .B(_4531__bF_buf3), .Y(_2822_) );
AOI22X1 AOI22X1_150 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_21_), .C(instr_rdcycleh_bF_buf0), .D(count_cycle_53_), .Y(_2823_) );
OAI21X1 OAI21X1_3421 ( .A(_4529_), .B(_1305_), .C(_2823_), .Y(_2824_) );
OAI21X1 OAI21X1_3422 ( .A(_2822_), .B(_2824_), .C(cpu_state_2_bF_buf2_), .Y(_2825_) );
OAI21X1 OAI21X1_3423 ( .A(_4575__bF_buf2), .B(_5217_), .C(_2825_), .Y(_2826_) );
AOI21X1 AOI21X1_963 ( .A(_4447__bF_buf3), .B(_2821_), .C(_2826_), .Y(_2827_) );
OAI21X1 OAI21X1_3424 ( .A(_2819_), .B(_2820_), .C(_2827_), .Y(_83__21_) );
NOR2X1 NOR2X1_1321 ( .A(_2803_), .B(_2816_), .Y(_2828_) );
INVX1 INVX1_1232 ( .A(_2828_), .Y(_2829_) );
AOI21X1 AOI21X1_964 ( .A(_2801_), .B(_2815_), .C(_2814_), .Y(_2830_) );
OAI21X1 OAI21X1_3425 ( .A(_2799_), .B(_2829_), .C(_2830_), .Y(_2831_) );
NOR2X1 NOR2X1_1322 ( .A(reg_pc_22_), .B(decoded_imm_22_), .Y(_2832_) );
AND2X2 AND2X2_214 ( .A(reg_pc_22_), .B(decoded_imm_22_), .Y(_2833_) );
NOR2X1 NOR2X1_1323 ( .A(_2832_), .B(_2833_), .Y(_2834_) );
AND2X2 AND2X2_215 ( .A(_2831_), .B(_2834_), .Y(_2835_) );
OAI21X1 OAI21X1_3426 ( .A(_2831_), .B(_2834_), .C(cpu_state_3_bF_buf1_), .Y(_2836_) );
INVX1 INVX1_1233 ( .A(mem_rdata[22]), .Y(_2837_) );
OAI21X1 OAI21X1_3427 ( .A(_2837_), .B(_2753_), .C(_2754_), .Y(_2838_) );
AND2X2 AND2X2_216 ( .A(_2421_), .B(count_instr_54_), .Y(_2839_) );
NAND2X1 NAND2X1_1058 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_22_), .Y(_2840_) );
NAND2X1 NAND2X1_1059 ( .A(instr_rdcycleh_bF_buf3), .B(count_cycle_54_), .Y(_2841_) );
NAND2X1 NAND2X1_1060 ( .A(instr_rdinstr_bF_buf2), .B(count_instr_22_), .Y(_2842_) );
NAND3X1 NAND3X1_104 ( .A(_2840_), .B(_2841_), .C(_2842_), .Y(_2843_) );
OAI21X1 OAI21X1_3428 ( .A(_2839_), .B(_2843_), .C(cpu_state_2_bF_buf1_), .Y(_2844_) );
OAI21X1 OAI21X1_3429 ( .A(_4575__bF_buf1), .B(_9021_), .C(_2844_), .Y(_2845_) );
AOI21X1 AOI21X1_965 ( .A(_4447__bF_buf2), .B(_2838_), .C(_2845_), .Y(_2846_) );
OAI21X1 OAI21X1_3430 ( .A(_2835_), .B(_2836_), .C(_2846_), .Y(_83__22_) );
NOR2X1 NOR2X1_1324 ( .A(_2833_), .B(_2835_), .Y(_2847_) );
NOR2X1 NOR2X1_1325 ( .A(reg_pc_23_), .B(decoded_imm_23_), .Y(_2848_) );
NOR2X1 NOR2X1_1326 ( .A(_4826_), .B(_1659_), .Y(_2849_) );
NOR2X1 NOR2X1_1327 ( .A(_2848_), .B(_2849_), .Y(_2850_) );
INVX1 INVX1_1234 ( .A(_2850_), .Y(_2851_) );
AND2X2 AND2X2_217 ( .A(_2847_), .B(_2851_), .Y(_2852_) );
OAI21X1 OAI21X1_3431 ( .A(_2847_), .B(_2851_), .C(cpu_state_3_bF_buf0_), .Y(_2853_) );
OAI21X1 OAI21X1_3432 ( .A(_1513_), .B(_2753_), .C(_2754_), .Y(_2854_) );
INVX1 INVX1_1235 ( .A(count_cycle_55_), .Y(_2855_) );
NOR2X1 NOR2X1_1328 ( .A(_1735_), .B(_2855_), .Y(_2856_) );
AOI22X1 AOI22X1_151 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_23_), .C(instr_rdinstr_bF_buf1), .D(count_instr_23_), .Y(_2857_) );
OAI21X1 OAI21X1_3433 ( .A(_4531__bF_buf2), .B(_1461_), .C(_2857_), .Y(_2858_) );
OAI21X1 OAI21X1_3434 ( .A(_2858_), .B(_2856_), .C(cpu_state_2_bF_buf0_), .Y(_2859_) );
OAI21X1 OAI21X1_3435 ( .A(_4575__bF_buf0), .B(_9091_), .C(_2859_), .Y(_2860_) );
AOI21X1 AOI21X1_966 ( .A(_4447__bF_buf1), .B(_2854_), .C(_2860_), .Y(_2861_) );
OAI21X1 OAI21X1_3436 ( .A(_2852_), .B(_2853_), .C(_2861_), .Y(_83__23_) );
NAND2X1 NAND2X1_1061 ( .A(_2834_), .B(_2850_), .Y(_2862_) );
AOI21X1 AOI21X1_967 ( .A(_2833_), .B(_2850_), .C(_2849_), .Y(_2863_) );
OAI21X1 OAI21X1_3437 ( .A(_2830_), .B(_2862_), .C(_2863_), .Y(_2864_) );
NOR2X1 NOR2X1_1329 ( .A(_2862_), .B(_2829_), .Y(_2865_) );
AOI21X1 AOI21X1_968 ( .A(_2865_), .B(_2798_), .C(_2864_), .Y(_2866_) );
NAND2X1 NAND2X1_1062 ( .A(_2865_), .B(_2796_), .Y(_2867_) );
OAI21X1 OAI21X1_3438 ( .A(_2728_), .B(_2867_), .C(_2866_), .Y(_2868_) );
NAND2X1 NAND2X1_1063 ( .A(_4841_), .B(_9440_), .Y(_2869_) );
NOR2X1 NOR2X1_1330 ( .A(_4841_), .B(_9440_), .Y(_2870_) );
INVX1 INVX1_1236 ( .A(_2870_), .Y(_2871_) );
AND2X2 AND2X2_218 ( .A(_2871_), .B(_2869_), .Y(_2872_) );
NOR2X1 NOR2X1_1331 ( .A(_2872_), .B(_2868_), .Y(_2873_) );
INVX1 INVX1_1237 ( .A(_2867_), .Y(_2874_) );
OAI21X1 OAI21X1_3439 ( .A(_2721_), .B(_2719_), .C(_2874_), .Y(_2875_) );
AND2X2 AND2X2_219 ( .A(_2875_), .B(_2866_), .Y(_2876_) );
INVX1 INVX1_1238 ( .A(_2872_), .Y(_2877_) );
OAI21X1 OAI21X1_3440 ( .A(_2876_), .B(_2877_), .C(cpu_state_3_bF_buf4_), .Y(_2878_) );
OAI21X1 OAI21X1_3441 ( .A(_1529_), .B(_2753_), .C(_2754_), .Y(_2879_) );
NOR2X1 NOR2X1_1332 ( .A(_1465_), .B(_4531__bF_buf1), .Y(_2880_) );
AOI22X1 AOI22X1_152 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_24_), .C(instr_rdcycleh_bF_buf2), .D(count_cycle_56_), .Y(_2881_) );
OAI21X1 OAI21X1_3442 ( .A(_4529_), .B(_1317_), .C(_2881_), .Y(_2882_) );
OAI21X1 OAI21X1_3443 ( .A(_2880_), .B(_2882_), .C(cpu_state_2_bF_buf5_), .Y(_2883_) );
OAI21X1 OAI21X1_3444 ( .A(_4575__bF_buf4), .B(_5032_), .C(_2883_), .Y(_2884_) );
AOI21X1 AOI21X1_969 ( .A(_4447__bF_buf0), .B(_2879_), .C(_2884_), .Y(_2885_) );
OAI21X1 OAI21X1_3445 ( .A(_2878_), .B(_2873_), .C(_2885_), .Y(_83__24_) );
NOR2X1 NOR2X1_1333 ( .A(reg_pc_25_), .B(decoded_imm_25_), .Y(_2886_) );
NOR2X1 NOR2X1_1334 ( .A(_4877_), .B(_9520_), .Y(_2887_) );
NOR2X1 NOR2X1_1335 ( .A(_2886_), .B(_2887_), .Y(_2888_) );
INVX1 INVX1_1239 ( .A(_2888_), .Y(_2889_) );
NOR2X1 NOR2X1_1336 ( .A(_2889_), .B(_2877_), .Y(_2890_) );
INVX1 INVX1_1240 ( .A(_2890_), .Y(_2891_) );
NOR2X1 NOR2X1_1337 ( .A(_2891_), .B(_2876_), .Y(_2892_) );
OAI21X1 OAI21X1_3446 ( .A(_2876_), .B(_2877_), .C(_2871_), .Y(_2893_) );
NOR2X1 NOR2X1_1338 ( .A(_2871_), .B(_2889_), .Y(_2894_) );
NOR2X1 NOR2X1_1339 ( .A(_4555_), .B(_2894_), .Y(_2895_) );
OAI21X1 OAI21X1_3447 ( .A(_2893_), .B(_2888_), .C(_2895_), .Y(_2896_) );
OAI21X1 OAI21X1_3448 ( .A(_1516_), .B(_2753_), .C(_2754_), .Y(_2897_) );
NAND2X1 NAND2X1_1064 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_25_), .Y(_2898_) );
NAND2X1 NAND2X1_1065 ( .A(instr_rdcycleh_bF_buf1), .B(count_cycle_57_), .Y(_2899_) );
NAND2X1 NAND2X1_1066 ( .A(instr_rdinstr_bF_buf0), .B(count_instr_25_), .Y(_2900_) );
NAND3X1 NAND3X1_105 ( .A(_2898_), .B(_2899_), .C(_2900_), .Y(_2901_) );
AOI21X1 AOI21X1_970 ( .A(count_instr_57_), .B(_2421_), .C(_2901_), .Y(_2902_) );
OAI22X1 OAI22X1_284 ( .A(_4575__bF_buf3), .B(_5027_), .C(_2902_), .D(_4538__bF_buf2), .Y(_2903_) );
AOI21X1 AOI21X1_971 ( .A(_4447__bF_buf3), .B(_2897_), .C(_2903_), .Y(_2904_) );
OAI21X1 OAI21X1_3449 ( .A(_2896_), .B(_2892_), .C(_2904_), .Y(_83__25_) );
NOR2X1 NOR2X1_1340 ( .A(_2887_), .B(_2894_), .Y(_2905_) );
OAI21X1 OAI21X1_3450 ( .A(_2876_), .B(_2891_), .C(_2905_), .Y(_2906_) );
NAND2X1 NAND2X1_1067 ( .A(_4860_), .B(_9607_), .Y(_2907_) );
NOR2X1 NOR2X1_1341 ( .A(_4860_), .B(_9607_), .Y(_2908_) );
INVX1 INVX1_1241 ( .A(_2908_), .Y(_2909_) );
AND2X2 AND2X2_220 ( .A(_2909_), .B(_2907_), .Y(_2910_) );
NOR2X1 NOR2X1_1342 ( .A(_2910_), .B(_2906_), .Y(_2911_) );
INVX1 INVX1_1242 ( .A(_2906_), .Y(_2912_) );
INVX1 INVX1_1243 ( .A(_2910_), .Y(_2913_) );
OAI21X1 OAI21X1_3451 ( .A(_2912_), .B(_2913_), .C(cpu_state_3_bF_buf3_), .Y(_2914_) );
OAI21X1 OAI21X1_3452 ( .A(_1504_), .B(_2753_), .C(_2754_), .Y(_2915_) );
AND2X2 AND2X2_221 ( .A(_2421_), .B(count_instr_58_), .Y(_2916_) );
NAND2X1 NAND2X1_1068 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_26_), .Y(_2917_) );
NAND2X1 NAND2X1_1069 ( .A(instr_rdinstr_bF_buf4), .B(count_instr_26_), .Y(_2918_) );
NAND2X1 NAND2X1_1070 ( .A(instr_rdcycleh_bF_buf0), .B(count_cycle_58_), .Y(_2919_) );
NAND3X1 NAND3X1_106 ( .A(_2917_), .B(_2918_), .C(_2919_), .Y(_2920_) );
OAI21X1 OAI21X1_3453 ( .A(_2916_), .B(_2920_), .C(cpu_state_2_bF_buf4_), .Y(_2921_) );
OAI21X1 OAI21X1_3454 ( .A(_4575__bF_buf2), .B(_5021_), .C(_2921_), .Y(_2922_) );
AOI21X1 AOI21X1_972 ( .A(_4447__bF_buf2), .B(_2915_), .C(_2922_), .Y(_2923_) );
OAI21X1 OAI21X1_3455 ( .A(_2914_), .B(_2911_), .C(_2923_), .Y(_83__26_) );
XOR2X1 XOR2X1_11 ( .A(reg_pc_27_), .B(decoded_imm_27_), .Y(_2924_) );
OAI21X1 OAI21X1_3456 ( .A(_2912_), .B(_2913_), .C(_2909_), .Y(_2925_) );
NOR2X1 NOR2X1_1343 ( .A(_2924_), .B(_2925_), .Y(_2926_) );
INVX1 INVX1_1244 ( .A(_2924_), .Y(_2927_) );
NOR2X1 NOR2X1_1344 ( .A(_2927_), .B(_2913_), .Y(_2928_) );
INVX1 INVX1_1245 ( .A(_2928_), .Y(_2929_) );
NOR2X1 NOR2X1_1345 ( .A(_2909_), .B(_2927_), .Y(_2930_) );
NOR2X1 NOR2X1_1346 ( .A(_4555_), .B(_2930_), .Y(_2931_) );
OAI21X1 OAI21X1_3457 ( .A(_2912_), .B(_2929_), .C(_2931_), .Y(_2932_) );
OAI21X1 OAI21X1_3458 ( .A(_1501_), .B(_2753_), .C(_2754_), .Y(_2933_) );
AND2X2 AND2X2_222 ( .A(_2421_), .B(count_instr_59_), .Y(_2934_) );
INVX1 INVX1_1246 ( .A(count_cycle_59_), .Y(_2935_) );
AOI22X1 AOI22X1_153 ( .A(instr_rdcycle_bF_buf0), .B(count_cycle_27_), .C(instr_rdinstr_bF_buf3), .D(count_instr_27_), .Y(_2936_) );
OAI21X1 OAI21X1_3459 ( .A(_1735_), .B(_2935_), .C(_2936_), .Y(_2937_) );
OAI21X1 OAI21X1_3460 ( .A(_2934_), .B(_2937_), .C(cpu_state_2_bF_buf3_), .Y(_2938_) );
OAI21X1 OAI21X1_3461 ( .A(_4575__bF_buf1), .B(_5016_), .C(_2938_), .Y(_2939_) );
AOI21X1 AOI21X1_973 ( .A(_4447__bF_buf1), .B(_2933_), .C(_2939_), .Y(_2940_) );
OAI21X1 OAI21X1_3462 ( .A(_2926_), .B(_2932_), .C(_2940_), .Y(_83__27_) );
AOI21X1 AOI21X1_974 ( .A(reg_pc_27_), .B(decoded_imm_27_), .C(_2930_), .Y(_2941_) );
OAI21X1 OAI21X1_3463 ( .A(_2929_), .B(_2905_), .C(_2941_), .Y(_2942_) );
NOR2X1 NOR2X1_1347 ( .A(_2929_), .B(_2891_), .Y(_2943_) );
AOI21X1 AOI21X1_975 ( .A(_2943_), .B(_2868_), .C(_2942_), .Y(_2944_) );
NOR2X1 NOR2X1_1348 ( .A(reg_pc_28_), .B(decoded_imm_28_), .Y(_2945_) );
NOR2X1 NOR2X1_1349 ( .A(_1215_), .B(_9770_), .Y(_2946_) );
OAI21X1 OAI21X1_3464 ( .A(_2945_), .B(_2946_), .C(_2944_), .Y(_2947_) );
NOR2X1 NOR2X1_1350 ( .A(_2945_), .B(_2946_), .Y(_2948_) );
INVX1 INVX1_1247 ( .A(_2948_), .Y(_2949_) );
OR2X2 OR2X2_44 ( .A(_2944_), .B(_2949_), .Y(_2950_) );
NAND2X1 NAND2X1_1071 ( .A(_2947_), .B(_2950_), .Y(_2951_) );
OAI21X1 OAI21X1_3465 ( .A(_1519_), .B(_2753_), .C(_2754_), .Y(_2952_) );
INVX1 INVX1_1248 ( .A(count_cycle_60_), .Y(_2953_) );
NOR2X1 NOR2X1_1351 ( .A(_1735_), .B(_2953_), .Y(_2954_) );
AOI22X1 AOI22X1_154 ( .A(instr_rdcycle_bF_buf4), .B(count_cycle_28_), .C(instr_rdinstr_bF_buf2), .D(count_instr_28_), .Y(_2955_) );
OAI21X1 OAI21X1_3466 ( .A(_4531__bF_buf0), .B(_1479_), .C(_2955_), .Y(_2956_) );
OAI21X1 OAI21X1_3467 ( .A(_2956_), .B(_2954_), .C(cpu_state_2_bF_buf2_), .Y(_2957_) );
OAI21X1 OAI21X1_3468 ( .A(_4575__bF_buf0), .B(_5004_), .C(_2957_), .Y(_2958_) );
AOI21X1 AOI21X1_976 ( .A(_4447__bF_buf0), .B(_2952_), .C(_2958_), .Y(_2959_) );
OAI21X1 OAI21X1_3469 ( .A(_2951_), .B(_4555_), .C(_2959_), .Y(_83__28_) );
OAI21X1 OAI21X1_3470 ( .A(_1215_), .B(_9770_), .C(_2950_), .Y(_2960_) );
NOR2X1 NOR2X1_1352 ( .A(reg_pc_29_), .B(decoded_imm_29_), .Y(_2961_) );
NOR2X1 NOR2X1_1353 ( .A(_4890_), .B(_9859_), .Y(_2962_) );
NOR2X1 NOR2X1_1354 ( .A(_2961_), .B(_2962_), .Y(_2963_) );
AND2X2 AND2X2_223 ( .A(_2960_), .B(_2963_), .Y(_2964_) );
OAI21X1 OAI21X1_3471 ( .A(_2960_), .B(_2963_), .C(cpu_state_3_bF_buf2_), .Y(_2965_) );
OAI21X1 OAI21X1_3472 ( .A(_1522_), .B(_2753_), .C(_2754_), .Y(_2966_) );
INVX1 INVX1_1249 ( .A(count_cycle_61_), .Y(_2967_) );
NOR2X1 NOR2X1_1355 ( .A(_1735_), .B(_2967_), .Y(_2968_) );
AOI22X1 AOI22X1_155 ( .A(instr_rdcycle_bF_buf3), .B(count_cycle_29_), .C(instr_rdinstr_bF_buf1), .D(count_instr_29_), .Y(_2969_) );
OAI21X1 OAI21X1_3473 ( .A(_4531__bF_buf4), .B(_1482_), .C(_2969_), .Y(_2970_) );
OAI21X1 OAI21X1_3474 ( .A(_2970_), .B(_2968_), .C(cpu_state_2_bF_buf1_), .Y(_2971_) );
OAI21X1 OAI21X1_3475 ( .A(_4575__bF_buf4), .B(_5009_), .C(_2971_), .Y(_2972_) );
AOI21X1 AOI21X1_977 ( .A(_4447__bF_buf3), .B(_2966_), .C(_2972_), .Y(_2973_) );
OAI21X1 OAI21X1_3476 ( .A(_2964_), .B(_2965_), .C(_2973_), .Y(_83__29_) );
AOI21X1 AOI21X1_978 ( .A(_2946_), .B(_2963_), .C(_2962_), .Y(_2974_) );
NAND2X1 NAND2X1_1072 ( .A(_2948_), .B(_2963_), .Y(_2975_) );
OAI21X1 OAI21X1_3477 ( .A(_2944_), .B(_2975_), .C(_2974_), .Y(_2976_) );
NOR2X1 NOR2X1_1356 ( .A(_4898_), .B(_9943_), .Y(_2977_) );
NOR2X1 NOR2X1_1357 ( .A(reg_pc_30_), .B(decoded_imm_30_), .Y(_2978_) );
NOR2X1 NOR2X1_1358 ( .A(_2978_), .B(_2977_), .Y(_2979_) );
AND2X2 AND2X2_224 ( .A(_2976_), .B(_2979_), .Y(_2980_) );
OAI21X1 OAI21X1_3478 ( .A(_2976_), .B(_2979_), .C(cpu_state_3_bF_buf1_), .Y(_2981_) );
OAI21X1 OAI21X1_3479 ( .A(_1498_), .B(_2753_), .C(_2754_), .Y(_2982_) );
INVX1 INVX1_1250 ( .A(count_cycle_62_), .Y(_2983_) );
NOR2X1 NOR2X1_1359 ( .A(_1735_), .B(_2983_), .Y(_2984_) );
AOI22X1 AOI22X1_156 ( .A(instr_rdcycle_bF_buf2), .B(count_cycle_30_), .C(instr_rdinstr_bF_buf0), .D(count_instr_30_), .Y(_2985_) );
OAI21X1 OAI21X1_3480 ( .A(_4531__bF_buf3), .B(_1489_), .C(_2985_), .Y(_2986_) );
OAI21X1 OAI21X1_3481 ( .A(_2986_), .B(_2984_), .C(cpu_state_2_bF_buf0_), .Y(_2987_) );
OAI21X1 OAI21X1_3482 ( .A(_4575__bF_buf3), .B(_4998_), .C(_2987_), .Y(_2988_) );
AOI21X1 AOI21X1_979 ( .A(_4447__bF_buf2), .B(_2982_), .C(_2988_), .Y(_2989_) );
OAI21X1 OAI21X1_3483 ( .A(_2980_), .B(_2981_), .C(_2989_), .Y(_83__30_) );
AOI21X1 AOI21X1_980 ( .A(_2979_), .B(_2976_), .C(_2977_), .Y(_2990_) );
XOR2X1 XOR2X1_12 ( .A(reg_pc_31_), .B(decoded_imm_31_), .Y(_2991_) );
INVX1 INVX1_1251 ( .A(_2991_), .Y(_2992_) );
AND2X2 AND2X2_225 ( .A(_2990_), .B(_2992_), .Y(_2993_) );
OAI21X1 OAI21X1_3484 ( .A(_2990_), .B(_2992_), .C(cpu_state_3_bF_buf0_), .Y(_2994_) );
OAI21X1 OAI21X1_3485 ( .A(_1525_), .B(_2753_), .C(_2754_), .Y(_2995_) );
AND2X2 AND2X2_226 ( .A(_2421_), .B(count_instr_63_), .Y(_2996_) );
AOI22X1 AOI22X1_157 ( .A(instr_rdcycle_bF_buf1), .B(count_cycle_31_), .C(instr_rdcycleh_bF_buf3), .D(count_cycle_63_), .Y(_2997_) );
OAI21X1 OAI21X1_3486 ( .A(_4529_), .B(_1350_), .C(_2997_), .Y(_2998_) );
OAI21X1 OAI21X1_3487 ( .A(_2996_), .B(_2998_), .C(cpu_state_2_bF_buf5_), .Y(_2999_) );
OAI21X1 OAI21X1_3488 ( .A(_4575__bF_buf2), .B(_4991_), .C(_2999_), .Y(_3000_) );
AOI21X1 AOI21X1_981 ( .A(_4447__bF_buf1), .B(_2995_), .C(_3000_), .Y(_3001_) );
OAI21X1 OAI21X1_3489 ( .A(_2993_), .B(_2994_), .C(_3001_), .Y(_83__31_) );
INVX1 INVX1_1252 ( .A(is_compare), .Y(_3002_) );
INVX1 INVX1_1253 ( .A(_5255_), .Y(_3003_) );
NAND2X1 NAND2X1_1073 ( .A(_5253_), .B(_3003_), .Y(_3004_) );
NOR2X1 NOR2X1_1360 ( .A(instr_ori), .B(instr_or), .Y(_3005_) );
INVX1 INVX1_1254 ( .A(_3005__bF_buf4), .Y(_3006_) );
NOR2X1 NOR2X1_1361 ( .A(instr_andi), .B(instr_and), .Y(_3007_) );
INVX1 INVX1_1255 ( .A(_3007__bF_buf4), .Y(_3008_) );
AOI22X1 AOI22X1_158 ( .A(_3008_), .B(_5254_), .C(_3003_), .D(_3006_), .Y(_3009_) );
NOR2X1 NOR2X1_1362 ( .A(instr_xori), .B(instr_xor), .Y(_3010_) );
INVX1 INVX1_1256 ( .A(_3010_), .Y(_3011_) );
NOR2X1 NOR2X1_1363 ( .A(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .B(_3011__bF_buf4), .Y(_3012_) );
OAI21X1 OAI21X1_3490 ( .A(_3012_), .B(_3004_), .C(_3009_), .Y(_3013_) );
NAND2X1 NAND2X1_1074 ( .A(_10734__15_), .B(_10728__0_bF_buf3_), .Y(_3014_) );
OAI21X1 OAI21X1_3491 ( .A(_5203_), .B(_10728__0_bF_buf2_), .C(_3014_), .Y(_3015_) );
NAND2X1 NAND2X1_1075 ( .A(_10734__13_), .B(_10728__0_bF_buf1_), .Y(_3016_) );
OAI21X1 OAI21X1_3492 ( .A(_5197_), .B(_10728__0_bF_buf0_), .C(_3016_), .Y(_3017_) );
MUX2X1 MUX2X1_261 ( .A(_3017_), .B(_3015_), .S(_5140__bF_buf0), .Y(_3018_) );
NAND2X1 NAND2X1_1076 ( .A(_10734__11_), .B(_10728__0_bF_buf7_), .Y(_3019_) );
OAI21X1 OAI21X1_3493 ( .A(_5121_), .B(_10728__0_bF_buf6_), .C(_3019_), .Y(_3020_) );
NAND2X1 NAND2X1_1077 ( .A(_10734__9_), .B(_10728__0_bF_buf5_), .Y(_3021_) );
OAI21X1 OAI21X1_3494 ( .A(_5187_), .B(_10728__0_bF_buf4_), .C(_3021_), .Y(_3022_) );
MUX2X1 MUX2X1_262 ( .A(_3022_), .B(_3020_), .S(_5140__bF_buf5), .Y(_3023_) );
MUX2X1 MUX2X1_263 ( .A(_3023_), .B(_3018_), .S(_5131__bF_buf0), .Y(_3024_) );
NOR2X1 NOR2X1_1364 ( .A(_5856__bF_buf1), .B(_3024_), .Y(_3025_) );
NAND2X1 NAND2X1_1078 ( .A(_10734__7_), .B(_10728__0_bF_buf3_), .Y(_3026_) );
OAI21X1 OAI21X1_3495 ( .A(_5174_), .B(_10728__0_bF_buf2_), .C(_3026_), .Y(_3027_) );
NAND2X1 NAND2X1_1079 ( .A(_10734__5_), .B(_10728__0_bF_buf1_), .Y(_3028_) );
OAI21X1 OAI21X1_3496 ( .A(_5180_), .B(_10728__0_bF_buf0_), .C(_3028_), .Y(_3029_) );
MUX2X1 MUX2X1_264 ( .A(_3029_), .B(_3027_), .S(_5140__bF_buf4), .Y(_3030_) );
NAND2X1 NAND2X1_1080 ( .A(_10734__3_), .B(_10728__0_bF_buf7_), .Y(_3031_) );
OAI21X1 OAI21X1_3497 ( .A(_5148_), .B(_10728__0_bF_buf6_), .C(_3031_), .Y(_3032_) );
AOI21X1 AOI21X1_982 ( .A(_4490_), .B(_10728__0_bF_buf5_), .C(_5255_), .Y(_3033_) );
MUX2X1 MUX2X1_265 ( .A(_3033_), .B(_3032_), .S(_5140__bF_buf3), .Y(_3034_) );
MUX2X1 MUX2X1_266 ( .A(_3034_), .B(_3030_), .S(_5131__bF_buf5), .Y(_3035_) );
NOR2X1 NOR2X1_1365 ( .A(_10728__3_bF_buf4_), .B(_3035_), .Y(_3036_) );
OAI21X1 OAI21X1_3498 ( .A(_3036_), .B(_3025_), .C(_5859__bF_buf0), .Y(_3037_) );
INVX1 INVX1_1257 ( .A(_3012_), .Y(_3038_) );
NAND3X1 NAND3X1_107 ( .A(_3002_), .B(_3005__bF_buf3), .C(_3007__bF_buf3), .Y(_3039_) );
NOR2X1 NOR2X1_1366 ( .A(_3039_), .B(_3038_), .Y(_3040_) );
INVX1 INVX1_1258 ( .A(_3040_), .Y(_3041_) );
NAND2X1 NAND2X1_1081 ( .A(_10734__27_), .B(_10728__0_bF_buf4_), .Y(_3042_) );
OAI21X1 OAI21X1_3499 ( .A(_5021_), .B(_10728__0_bF_buf3_), .C(_3042_), .Y(_3043_) );
NAND2X1 NAND2X1_1082 ( .A(_10734__25_), .B(_10728__0_bF_buf2_), .Y(_3044_) );
OAI21X1 OAI21X1_3500 ( .A(_5032_), .B(_10728__0_bF_buf1_), .C(_3044_), .Y(_3045_) );
INVX1 INVX1_1259 ( .A(_3045_), .Y(_3046_) );
NAND2X1 NAND2X1_1083 ( .A(_5140__bF_buf2), .B(_3046_), .Y(_3047_) );
OAI21X1 OAI21X1_3501 ( .A(_5140__bF_buf1), .B(_3043_), .C(_3047_), .Y(_3048_) );
NAND2X1 NAND2X1_1084 ( .A(_10734__29_), .B(_10728__0_bF_buf0_), .Y(_3049_) );
OAI21X1 OAI21X1_3502 ( .A(_5004_), .B(_10728__0_bF_buf7_), .C(_3049_), .Y(_3050_) );
INVX1 INVX1_1260 ( .A(_3050_), .Y(_3051_) );
NAND2X1 NAND2X1_1085 ( .A(_10734__31_), .B(_10728__0_bF_buf6_), .Y(_3052_) );
OAI21X1 OAI21X1_3503 ( .A(_4998_), .B(_10728__0_bF_buf5_), .C(_3052_), .Y(_3053_) );
NAND2X1 NAND2X1_1086 ( .A(_10728__1_bF_buf0_), .B(_3053_), .Y(_3054_) );
OAI21X1 OAI21X1_3504 ( .A(_3051_), .B(_10728__1_bF_buf3_), .C(_3054_), .Y(_3055_) );
NAND2X1 NAND2X1_1087 ( .A(_10728__2_bF_buf1_), .B(_3055_), .Y(_3056_) );
OAI21X1 OAI21X1_3505 ( .A(_3048_), .B(_10728__2_bF_buf0_), .C(_3056_), .Y(_3057_) );
INVX1 INVX1_1261 ( .A(_3057_), .Y(_3058_) );
NAND2X1 NAND2X1_1088 ( .A(_10728__3_bF_buf3_), .B(_3058_), .Y(_3059_) );
NAND2X1 NAND2X1_1089 ( .A(_10734__23_), .B(_10728__0_bF_buf4_), .Y(_3060_) );
OAI21X1 OAI21X1_3506 ( .A(_9021_), .B(_10728__0_bF_buf3_), .C(_3060_), .Y(_3061_) );
NAND2X1 NAND2X1_1090 ( .A(_10734__21_), .B(_10728__0_bF_buf2_), .Y(_3062_) );
OAI21X1 OAI21X1_3507 ( .A(_5218_), .B(_10728__0_bF_buf1_), .C(_3062_), .Y(_3063_) );
INVX1 INVX1_1262 ( .A(_3063_), .Y(_3064_) );
NAND2X1 NAND2X1_1091 ( .A(_5140__bF_buf0), .B(_3064_), .Y(_3065_) );
OAI21X1 OAI21X1_3508 ( .A(_5140__bF_buf5), .B(_3061_), .C(_3065_), .Y(_3066_) );
NAND2X1 NAND2X1_1092 ( .A(_10734__19_), .B(_10728__0_bF_buf0_), .Y(_3067_) );
OAI21X1 OAI21X1_3509 ( .A(_5045_), .B(_10728__0_bF_buf7_), .C(_3067_), .Y(_3068_) );
NAND2X1 NAND2X1_1093 ( .A(_10734__17_), .B(_10728__0_bF_buf6_), .Y(_3069_) );
OAI21X1 OAI21X1_3510 ( .A(_5051_), .B(_10728__0_bF_buf5_), .C(_3069_), .Y(_3070_) );
MUX2X1 MUX2X1_267 ( .A(_3070_), .B(_3068_), .S(_5140__bF_buf4), .Y(_3071_) );
MUX2X1 MUX2X1_268 ( .A(_3066_), .B(_3071_), .S(_10728__2_bF_buf4_), .Y(_3072_) );
OAI21X1 OAI21X1_3511 ( .A(_10728__3_bF_buf2_), .B(_3072_), .C(_3059_), .Y(_3073_) );
AOI21X1 AOI21X1_983 ( .A(_10728__4_bF_buf4_), .B(_3073_), .C(_3041_), .Y(_3074_) );
AOI21X1 AOI21X1_984 ( .A(_3037_), .B(_3074_), .C(_3013_), .Y(_3075_) );
OAI21X1 OAI21X1_3512 ( .A(_5266_), .B(_3002_), .C(_3075_), .Y(alu_out_0_) );
NAND2X1 NAND2X1_1094 ( .A(_10734__30_), .B(_10728__0_bF_buf4_), .Y(_3076_) );
OAI21X1 OAI21X1_3513 ( .A(_5009_), .B(_10728__0_bF_buf3_), .C(_3076_), .Y(_3077_) );
NOR2X1 NOR2X1_1367 ( .A(_10728__0_bF_buf2_), .B(_4991_), .Y(_3078_) );
OAI21X1 OAI21X1_3514 ( .A(instr_srai), .B(instr_sra), .C(_10734__31_), .Y(_3079_) );
NAND2X1 NAND2X1_1095 ( .A(_10728__1_bF_buf2_), .B(_3079_), .Y(_3080_) );
OAI22X1 OAI22X1_285 ( .A(_10728__1_bF_buf1_), .B(_3077_), .C(_3080_), .D(_3078_), .Y(_3081_) );
NAND2X1 NAND2X1_1096 ( .A(_10734__28_), .B(_10728__0_bF_buf1_), .Y(_3082_) );
OAI21X1 OAI21X1_3515 ( .A(_5016_), .B(_10728__0_bF_buf0_), .C(_3082_), .Y(_3083_) );
INVX1 INVX1_1263 ( .A(_3083_), .Y(_3084_) );
NAND2X1 NAND2X1_1097 ( .A(_10734__26_), .B(_10728__0_bF_buf7_), .Y(_3085_) );
OAI21X1 OAI21X1_3516 ( .A(_5027_), .B(_10728__0_bF_buf6_), .C(_3085_), .Y(_3086_) );
NAND2X1 NAND2X1_1098 ( .A(_5140__bF_buf3), .B(_3086_), .Y(_3087_) );
OAI21X1 OAI21X1_3517 ( .A(_3084_), .B(_5140__bF_buf2), .C(_3087_), .Y(_3088_) );
NAND2X1 NAND2X1_1099 ( .A(_5131__bF_buf4), .B(_3088_), .Y(_3089_) );
OAI21X1 OAI21X1_3518 ( .A(_5131__bF_buf3), .B(_3081_), .C(_3089_), .Y(_3090_) );
INVX1 INVX1_1264 ( .A(_3090_), .Y(_3091_) );
NAND2X1 NAND2X1_1100 ( .A(_10734__20_), .B(_10728__0_bF_buf5_), .Y(_3092_) );
OAI21X1 OAI21X1_3519 ( .A(_5040_), .B(_10728__0_bF_buf4_), .C(_3092_), .Y(_3093_) );
NAND2X1 NAND2X1_1101 ( .A(_10734__18_), .B(_10728__0_bF_buf3_), .Y(_3094_) );
OAI21X1 OAI21X1_3520 ( .A(_5057_), .B(_10728__0_bF_buf2_), .C(_3094_), .Y(_3095_) );
INVX1 INVX1_1265 ( .A(_3095_), .Y(_3096_) );
NAND2X1 NAND2X1_1102 ( .A(_5140__bF_buf1), .B(_3096_), .Y(_3097_) );
OAI21X1 OAI21X1_3521 ( .A(_5140__bF_buf0), .B(_3093_), .C(_3097_), .Y(_3098_) );
NAND2X1 NAND2X1_1103 ( .A(_10734__22_), .B(_10728__0_bF_buf1_), .Y(_3099_) );
OAI21X1 OAI21X1_3522 ( .A(_5217_), .B(_10728__0_bF_buf0_), .C(_3099_), .Y(_3100_) );
INVX1 INVX1_1266 ( .A(_3100_), .Y(_3101_) );
NAND2X1 NAND2X1_1104 ( .A(_10734__24_), .B(_10728__0_bF_buf7_), .Y(_3102_) );
OAI21X1 OAI21X1_3523 ( .A(_9091_), .B(_10728__0_bF_buf6_), .C(_3102_), .Y(_3103_) );
NAND2X1 NAND2X1_1105 ( .A(_10728__1_bF_buf0_), .B(_3103_), .Y(_3104_) );
OAI21X1 OAI21X1_3524 ( .A(_3101_), .B(_10728__1_bF_buf3_), .C(_3104_), .Y(_3105_) );
NAND2X1 NAND2X1_1106 ( .A(_10728__2_bF_buf3_), .B(_3105_), .Y(_3106_) );
OAI21X1 OAI21X1_3525 ( .A(_3098_), .B(_10728__2_bF_buf2_), .C(_3106_), .Y(_3107_) );
NAND2X1 NAND2X1_1107 ( .A(_5856__bF_buf0), .B(_3107_), .Y(_3108_) );
OAI21X1 OAI21X1_3526 ( .A(_3091_), .B(_5856__bF_buf4), .C(_3108_), .Y(_3109_) );
NOR2X1 NOR2X1_1368 ( .A(_5859__bF_buf4), .B(_3109_), .Y(_3110_) );
NAND2X1 NAND2X1_1108 ( .A(_10734__16_), .B(_10728__0_bF_buf5_), .Y(_3111_) );
OAI21X1 OAI21X1_3527 ( .A(_5087_), .B(_10728__0_bF_buf4_), .C(_3111_), .Y(_3112_) );
INVX1 INVX1_1267 ( .A(_3112_), .Y(_3113_) );
NAND2X1 NAND2X1_1109 ( .A(_10734__14_), .B(_10728__0_bF_buf3_), .Y(_3114_) );
OAI21X1 OAI21X1_3528 ( .A(_5196_), .B(_10728__0_bF_buf2_), .C(_3114_), .Y(_3115_) );
NAND2X1 NAND2X1_1110 ( .A(_5140__bF_buf5), .B(_3115_), .Y(_3116_) );
OAI21X1 OAI21X1_3529 ( .A(_3113_), .B(_5140__bF_buf4), .C(_3116_), .Y(_3117_) );
NAND2X1 NAND2X1_1111 ( .A(_10734__12_), .B(_10728__0_bF_buf1_), .Y(_3118_) );
OAI21X1 OAI21X1_3530 ( .A(_5117_), .B(_10728__0_bF_buf0_), .C(_3118_), .Y(_3119_) );
INVX1 INVX1_1268 ( .A(_3119_), .Y(_3120_) );
NAND2X1 NAND2X1_1112 ( .A(_10734__10_), .B(_10728__0_bF_buf7_), .Y(_3121_) );
OAI21X1 OAI21X1_3531 ( .A(_5107_), .B(_10728__0_bF_buf6_), .C(_3121_), .Y(_3122_) );
NAND2X1 NAND2X1_1113 ( .A(_5140__bF_buf3), .B(_3122_), .Y(_3123_) );
OAI21X1 OAI21X1_3532 ( .A(_3120_), .B(_5140__bF_buf2), .C(_3123_), .Y(_3124_) );
INVX1 INVX1_1269 ( .A(_3124_), .Y(_3125_) );
NAND2X1 NAND2X1_1114 ( .A(_5131__bF_buf2), .B(_3125_), .Y(_3126_) );
OAI21X1 OAI21X1_3533 ( .A(_5131__bF_buf1), .B(_3117_), .C(_3126_), .Y(_3127_) );
NAND2X1 NAND2X1_1115 ( .A(_10734__4_), .B(_10728__0_bF_buf5_), .Y(_3128_) );
OAI21X1 OAI21X1_3534 ( .A(_5130_), .B(_10728__0_bF_buf4_), .C(_3128_), .Y(_3129_) );
INVX1 INVX1_1270 ( .A(_3129_), .Y(_3130_) );
NAND2X1 NAND2X1_1116 ( .A(_10734__2_), .B(_10728__0_bF_buf3_), .Y(_3131_) );
OAI21X1 OAI21X1_3535 ( .A(_4490_), .B(_10728__0_bF_buf2_), .C(_3131_), .Y(_3132_) );
AOI21X1 AOI21X1_985 ( .A(_5140__bF_buf1), .B(_3132_), .C(_10728__2_bF_buf1_), .Y(_3133_) );
OAI21X1 OAI21X1_3536 ( .A(_5140__bF_buf0), .B(_3130_), .C(_3133_), .Y(_3134_) );
NAND2X1 NAND2X1_1117 ( .A(_10734__8_), .B(_10728__0_bF_buf1_), .Y(_3135_) );
OAI21X1 OAI21X1_3537 ( .A(_5173_), .B(_10728__0_bF_buf0_), .C(_3135_), .Y(_3136_) );
INVX1 INVX1_1271 ( .A(_3136_), .Y(_3137_) );
NAND2X1 NAND2X1_1118 ( .A(_10734__6_), .B(_10728__0_bF_buf7_), .Y(_3138_) );
OAI21X1 OAI21X1_3538 ( .A(_5179_), .B(_10728__0_bF_buf6_), .C(_3138_), .Y(_3139_) );
NAND2X1 NAND2X1_1119 ( .A(_5140__bF_buf5), .B(_3139_), .Y(_3140_) );
OAI21X1 OAI21X1_3539 ( .A(_3137_), .B(_5140__bF_buf4), .C(_3140_), .Y(_3141_) );
OAI21X1 OAI21X1_3540 ( .A(_3141_), .B(_5131__bF_buf0), .C(_3134_), .Y(_3142_) );
MUX2X1 MUX2X1_269 ( .A(_3127_), .B(_3142_), .S(_10728__3_bF_buf1_), .Y(_3143_) );
OAI21X1 OAI21X1_3541 ( .A(_3143_), .B(_10728__4_bF_buf3_), .C(_3040_), .Y(_3144_) );
NAND3X1 NAND3X1_108 ( .A(instr_sub_bF_buf3), .B(_10728__0_bF_buf5_), .C(_4491_), .Y(_3145_) );
OAI21X1 OAI21X1_3542 ( .A(instr_sub_bF_buf2), .B(_5253_), .C(_3145_), .Y(_3146_) );
XNOR2X1 XNOR2X1_57 ( .A(_3146_), .B(_5145_), .Y(_3147_) );
NOR2X1 NOR2X1_1369 ( .A(_3010_), .B(_5145_), .Y(_3148_) );
OAI21X1 OAI21X1_3543 ( .A(instr_ori), .B(instr_or), .C(_5144_), .Y(_3149_) );
OAI21X1 OAI21X1_3544 ( .A(_5143_), .B(_3007__bF_buf2), .C(_3149_), .Y(_3150_) );
OR2X2 OR2X2_45 ( .A(_3148_), .B(_3150_), .Y(_3151_) );
AOI21X1 AOI21X1_986 ( .A(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3), .B(_3147_), .C(_3151_), .Y(_3152_) );
OAI21X1 OAI21X1_3545 ( .A(_3144_), .B(_3110_), .C(_3152_), .Y(alu_out_1_) );
MUX2X1 MUX2X1_270 ( .A(_3032_), .B(_3029_), .S(_5140__bF_buf3), .Y(_3153_) );
MUX2X1 MUX2X1_271 ( .A(_3027_), .B(_3022_), .S(_5140__bF_buf2), .Y(_3154_) );
MUX2X1 MUX2X1_272 ( .A(_3154_), .B(_3153_), .S(_10728__2_bF_buf0_), .Y(_3155_) );
NOR2X1 NOR2X1_1370 ( .A(_10728__3_bF_buf0_), .B(_3155_), .Y(_3156_) );
MUX2X1 MUX2X1_273 ( .A(_3070_), .B(_3015_), .S(_10728__1_bF_buf2_), .Y(_3157_) );
MUX2X1 MUX2X1_274 ( .A(_3020_), .B(_3017_), .S(_5140__bF_buf1), .Y(_3158_) );
MUX2X1 MUX2X1_275 ( .A(_3158_), .B(_3157_), .S(_5131__bF_buf5), .Y(_3159_) );
OAI21X1 OAI21X1_3546 ( .A(_3159_), .B(_5856__bF_buf3), .C(_5859__bF_buf3), .Y(_3160_) );
OAI21X1 OAI21X1_3547 ( .A(_3053_), .B(_10728__1_bF_buf1_), .C(_3080_), .Y(_3161_) );
NAND2X1 NAND2X1_1120 ( .A(_5140__bF_buf0), .B(_3043_), .Y(_3162_) );
OAI21X1 OAI21X1_3548 ( .A(_3051_), .B(_5140__bF_buf5), .C(_3162_), .Y(_3163_) );
NAND2X1 NAND2X1_1121 ( .A(_5131__bF_buf4), .B(_3163_), .Y(_3164_) );
OAI21X1 OAI21X1_3549 ( .A(_5131__bF_buf3), .B(_3161_), .C(_3164_), .Y(_3165_) );
INVX1 INVX1_1272 ( .A(_3165_), .Y(_3166_) );
NAND2X1 NAND2X1_1122 ( .A(_5140__bF_buf4), .B(_3061_), .Y(_3167_) );
OAI21X1 OAI21X1_3550 ( .A(_3046_), .B(_5140__bF_buf3), .C(_3167_), .Y(_3168_) );
INVX1 INVX1_1273 ( .A(_3168_), .Y(_3169_) );
NAND2X1 NAND2X1_1123 ( .A(_5140__bF_buf2), .B(_3068_), .Y(_3170_) );
OAI21X1 OAI21X1_3551 ( .A(_3064_), .B(_5140__bF_buf1), .C(_3170_), .Y(_3171_) );
NAND2X1 NAND2X1_1124 ( .A(_5131__bF_buf2), .B(_3171_), .Y(_3172_) );
OAI21X1 OAI21X1_3552 ( .A(_3169_), .B(_5131__bF_buf1), .C(_3172_), .Y(_3173_) );
NAND2X1 NAND2X1_1125 ( .A(_5856__bF_buf2), .B(_3173_), .Y(_3174_) );
OAI21X1 OAI21X1_3553 ( .A(_3166_), .B(_5856__bF_buf1), .C(_3174_), .Y(_3175_) );
NAND2X1 NAND2X1_1126 ( .A(_10728__4_bF_buf2_), .B(_3175_), .Y(_3176_) );
OAI21X1 OAI21X1_3554 ( .A(_3156_), .B(_3160_), .C(_3176_), .Y(_3177_) );
NAND2X1 NAND2X1_1127 ( .A(_3040_), .B(_3177_), .Y(_3178_) );
NOR2X1 NOR2X1_1371 ( .A(_5150_), .B(_5149_), .Y(_3179_) );
NAND2X1 NAND2X1_1128 ( .A(instr_sub_bF_buf1), .B(_5147_), .Y(_3180_) );
OAI21X1 OAI21X1_3555 ( .A(_4490_), .B(_5140__bF_buf0), .C(_5253_), .Y(_3181_) );
OAI21X1 OAI21X1_3556 ( .A(_10734__1_), .B(_10728__1_bF_buf0_), .C(_3181_), .Y(_3182_) );
OAI21X1 OAI21X1_3557 ( .A(instr_sub_bF_buf0), .B(_3182_), .C(_3180_), .Y(_3183_) );
INVX1 INVX1_1274 ( .A(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2), .Y(_3184_) );
AOI21X1 AOI21X1_987 ( .A(_3179_), .B(_3183_), .C(_3184_), .Y(_3185_) );
OAI21X1 OAI21X1_3558 ( .A(_3179_), .B(_3183_), .C(_3185_), .Y(_3186_) );
INVX1 INVX1_1275 ( .A(_5149_), .Y(_3187_) );
OAI22X1 OAI22X1_286 ( .A(_5150_), .B(_3005__bF_buf2), .C(_3187_), .D(_3007__bF_buf1), .Y(_3188_) );
AOI21X1 AOI21X1_988 ( .A(_3011__bF_buf3), .B(_3179_), .C(_3188_), .Y(_3189_) );
NAND3X1 NAND3X1_109 ( .A(_3186_), .B(_3189_), .C(_3178_), .Y(alu_out_2_) );
NAND2X1 NAND2X1_1129 ( .A(_5140__bF_buf5), .B(_3084_), .Y(_3190_) );
OAI21X1 OAI21X1_3559 ( .A(_5140__bF_buf4), .B(_3077_), .C(_3190_), .Y(_3191_) );
NAND2X1 NAND2X1_1130 ( .A(_5140__bF_buf3), .B(_3078_), .Y(_3192_) );
INVX1 INVX1_1276 ( .A(_3079_), .Y(_3193_) );
NOR2X1 NOR2X1_1372 ( .A(_5131__bF_buf0), .B(_3193_), .Y(_3194_) );
AOI22X1 AOI22X1_159 ( .A(_3192_), .B(_3194_), .C(_3191_), .D(_5131__bF_buf5), .Y(_3195_) );
INVX1 INVX1_1277 ( .A(_3195_), .Y(_3196_) );
INVX1 INVX1_1278 ( .A(_3086_), .Y(_3197_) );
NAND2X1 NAND2X1_1131 ( .A(_5140__bF_buf2), .B(_3103_), .Y(_3198_) );
OAI21X1 OAI21X1_3560 ( .A(_3197_), .B(_5140__bF_buf1), .C(_3198_), .Y(_3199_) );
INVX1 INVX1_1279 ( .A(_3199_), .Y(_3200_) );
NAND2X1 NAND2X1_1132 ( .A(_5140__bF_buf0), .B(_3093_), .Y(_3201_) );
OAI21X1 OAI21X1_3561 ( .A(_3101_), .B(_5140__bF_buf5), .C(_3201_), .Y(_3202_) );
NAND2X1 NAND2X1_1133 ( .A(_5131__bF_buf4), .B(_3202_), .Y(_3203_) );
OAI21X1 OAI21X1_3562 ( .A(_3200_), .B(_5131__bF_buf3), .C(_3203_), .Y(_3204_) );
NAND2X1 NAND2X1_1134 ( .A(_5856__bF_buf0), .B(_3204_), .Y(_3205_) );
OAI21X1 OAI21X1_3563 ( .A(_3196_), .B(_5856__bF_buf4), .C(_3205_), .Y(_3206_) );
NOR2X1 NOR2X1_1373 ( .A(_10728__1_bF_buf3_), .B(_3129_), .Y(_3207_) );
OAI21X1 OAI21X1_3564 ( .A(_3139_), .B(_5140__bF_buf4), .C(_5131__bF_buf2), .Y(_3208_) );
NAND2X1 NAND2X1_1135 ( .A(_5140__bF_buf3), .B(_3137_), .Y(_3209_) );
OAI21X1 OAI21X1_3565 ( .A(_5140__bF_buf2), .B(_3122_), .C(_3209_), .Y(_3210_) );
OAI22X1 OAI22X1_287 ( .A(_3207_), .B(_3208_), .C(_3210_), .D(_5131__bF_buf1), .Y(_3211_) );
NOR2X1 NOR2X1_1374 ( .A(_10728__3_bF_buf4_), .B(_3211_), .Y(_3212_) );
NAND2X1 NAND2X1_1136 ( .A(_5140__bF_buf1), .B(_3112_), .Y(_3213_) );
OAI21X1 OAI21X1_3566 ( .A(_3096_), .B(_5140__bF_buf0), .C(_3213_), .Y(_3214_) );
INVX1 INVX1_1280 ( .A(_3214_), .Y(_3215_) );
NAND2X1 NAND2X1_1137 ( .A(_10728__1_bF_buf2_), .B(_3115_), .Y(_3216_) );
OAI21X1 OAI21X1_3567 ( .A(_3120_), .B(_10728__1_bF_buf1_), .C(_3216_), .Y(_3217_) );
NAND2X1 NAND2X1_1138 ( .A(_5131__bF_buf0), .B(_3217_), .Y(_3218_) );
OAI21X1 OAI21X1_3568 ( .A(_3215_), .B(_5131__bF_buf5), .C(_3218_), .Y(_3219_) );
NOR2X1 NOR2X1_1375 ( .A(_5856__bF_buf3), .B(_3219_), .Y(_3220_) );
OAI21X1 OAI21X1_3569 ( .A(_3220_), .B(_3212_), .C(_5859__bF_buf2), .Y(_3221_) );
OAI21X1 OAI21X1_3570 ( .A(_5859__bF_buf1), .B(_3206_), .C(_3221_), .Y(_3222_) );
INVX1 INVX1_1281 ( .A(instr_sub_bF_buf4), .Y(_3223_) );
OAI21X1 OAI21X1_3571 ( .A(_5147_), .B(_3179_), .C(_5132_), .Y(_3224_) );
OAI21X1 OAI21X1_3572 ( .A(_3182_), .B(_5150_), .C(_3187_), .Y(_3225_) );
NAND2X1 NAND2X1_1139 ( .A(_3223__bF_buf3), .B(_3225_), .Y(_3226_) );
OAI21X1 OAI21X1_3573 ( .A(_3224_), .B(_3223__bF_buf2), .C(_3226_), .Y(_3227_) );
AOI21X1 AOI21X1_989 ( .A(_5137_), .B(_3227_), .C(_3184_), .Y(_3228_) );
OAI21X1 OAI21X1_3574 ( .A(_5137_), .B(_3227_), .C(_3228_), .Y(_3229_) );
OAI22X1 OAI22X1_288 ( .A(_3007__bF_buf0), .B(_5133_), .C(_5134_), .D(_3005__bF_buf1), .Y(_3230_) );
AOI21X1 AOI21X1_990 ( .A(_3011__bF_buf2), .B(_5137_), .C(_3230_), .Y(_3231_) );
AND2X2 AND2X2_227 ( .A(_3229_), .B(_3231_), .Y(_3232_) );
OAI21X1 OAI21X1_3575 ( .A(_3041_), .B(_3222_), .C(_3232_), .Y(alu_out_3_) );
NOR2X1 NOR2X1_1376 ( .A(_5169_), .B(_5168_), .Y(_3233_) );
NOR2X1 NOR2X1_1377 ( .A(_5139_), .B(_5152_), .Y(_3234_) );
NAND2X1 NAND2X1_1140 ( .A(instr_sub_bF_buf3), .B(_3234_), .Y(_3235_) );
OAI21X1 OAI21X1_3576 ( .A(_10734__3_), .B(_10728__3_bF_buf3_), .C(_3225_), .Y(_3236_) );
OAI21X1 OAI21X1_3577 ( .A(_5130_), .B(_5856__bF_buf2), .C(_3236_), .Y(_3237_) );
INVX1 INVX1_1282 ( .A(_3237_), .Y(_3238_) );
OAI21X1 OAI21X1_3578 ( .A(instr_sub_bF_buf2), .B(_3238_), .C(_3235_), .Y(_3239_) );
AOI21X1 AOI21X1_991 ( .A(_3233_), .B(_3239_), .C(_3184_), .Y(_3240_) );
OAI21X1 OAI21X1_3579 ( .A(_3233_), .B(_3239_), .C(_3240_), .Y(_3241_) );
MUX2X1 MUX2X1_276 ( .A(_3030_), .B(_3023_), .S(_5131__bF_buf4), .Y(_3242_) );
MUX2X1 MUX2X1_277 ( .A(_3071_), .B(_3018_), .S(_10728__2_bF_buf4_), .Y(_3243_) );
MUX2X1 MUX2X1_278 ( .A(_3243_), .B(_3242_), .S(_10728__3_bF_buf2_), .Y(_3244_) );
INVX1 INVX1_1283 ( .A(_3194_), .Y(_3245_) );
OAI21X1 OAI21X1_3580 ( .A(_3055_), .B(_10728__2_bF_buf3_), .C(_3245_), .Y(_3246_) );
MUX2X1 MUX2X1_279 ( .A(_3066_), .B(_3048_), .S(_5131__bF_buf3), .Y(_3247_) );
NAND2X1 NAND2X1_1141 ( .A(_5856__bF_buf1), .B(_3247_), .Y(_3248_) );
OAI21X1 OAI21X1_3581 ( .A(_5856__bF_buf0), .B(_3246_), .C(_3248_), .Y(_3249_) );
NAND2X1 NAND2X1_1142 ( .A(_10728__4_bF_buf1_), .B(_3249_), .Y(_3250_) );
OAI21X1 OAI21X1_3582 ( .A(_10728__4_bF_buf0_), .B(_3244_), .C(_3250_), .Y(_3251_) );
NAND2X1 NAND2X1_1143 ( .A(_3040_), .B(_3251_), .Y(_3252_) );
OAI22X1 OAI22X1_289 ( .A(_3007__bF_buf4), .B(_5167_), .C(_5169_), .D(_3005__bF_buf0), .Y(_3253_) );
AOI21X1 AOI21X1_992 ( .A(_3011__bF_buf1), .B(_3233_), .C(_3253_), .Y(_3254_) );
NAND3X1 NAND3X1_110 ( .A(_3252_), .B(_3254_), .C(_3241_), .Y(alu_out_4_) );
NOR2X1 NOR2X1_1378 ( .A(_3233_), .B(_3234_), .Y(_3255_) );
OAI21X1 OAI21X1_3583 ( .A(_3255_), .B(_5181_), .C(instr_sub_bF_buf1), .Y(_3256_) );
INVX1 INVX1_1284 ( .A(_3233_), .Y(_3257_) );
OAI21X1 OAI21X1_3584 ( .A(_3238_), .B(_3257_), .C(_5167_), .Y(_3258_) );
OAI21X1 OAI21X1_3585 ( .A(instr_sub_bF_buf0), .B(_3258_), .C(_3256_), .Y(_3259_) );
AND2X2 AND2X2_228 ( .A(_3259_), .B(_5166_), .Y(_3260_) );
OAI21X1 OAI21X1_3586 ( .A(_3259_), .B(_5166_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1), .Y(_3261_) );
NAND2X1 NAND2X1_1144 ( .A(_10728__2_bF_buf2_), .B(_3193_), .Y(_3262_) );
OAI21X1 OAI21X1_3587 ( .A(_3081_), .B(_10728__2_bF_buf1_), .C(_3262_), .Y(_3263_) );
INVX1 INVX1_1285 ( .A(_3263_), .Y(_3264_) );
INVX1 INVX1_1286 ( .A(_3088_), .Y(_3265_) );
NAND2X1 NAND2X1_1145 ( .A(_5131__bF_buf2), .B(_3105_), .Y(_3266_) );
OAI21X1 OAI21X1_3588 ( .A(_3265_), .B(_5131__bF_buf1), .C(_3266_), .Y(_3267_) );
NAND2X1 NAND2X1_1146 ( .A(_5856__bF_buf4), .B(_3267_), .Y(_3268_) );
OAI21X1 OAI21X1_3589 ( .A(_3264_), .B(_5856__bF_buf3), .C(_3268_), .Y(_3269_) );
NAND2X1 NAND2X1_1147 ( .A(_5131__bF_buf0), .B(_3117_), .Y(_3270_) );
OAI21X1 OAI21X1_3590 ( .A(_3098_), .B(_5131__bF_buf5), .C(_3270_), .Y(_3271_) );
NAND2X1 NAND2X1_1148 ( .A(_5131__bF_buf4), .B(_3141_), .Y(_3272_) );
OAI21X1 OAI21X1_3591 ( .A(_3125_), .B(_5131__bF_buf3), .C(_3272_), .Y(_3273_) );
MUX2X1 MUX2X1_280 ( .A(_3273_), .B(_3271_), .S(_5856__bF_buf2), .Y(_3274_) );
AOI21X1 AOI21X1_993 ( .A(_5859__bF_buf0), .B(_3274_), .C(_3041_), .Y(_3275_) );
OAI21X1 OAI21X1_3592 ( .A(_5859__bF_buf4), .B(_3269_), .C(_3275_), .Y(_3276_) );
OAI22X1 OAI22X1_290 ( .A(_3007__bF_buf3), .B(_5163_), .C(_5162_), .D(_3005__bF_buf4), .Y(_3277_) );
AOI21X1 AOI21X1_994 ( .A(_3011__bF_buf0), .B(_5165_), .C(_3277_), .Y(_3278_) );
AND2X2 AND2X2_229 ( .A(_3276_), .B(_3278_), .Y(_3279_) );
OAI21X1 OAI21X1_3593 ( .A(_3260_), .B(_3261_), .C(_3279_), .Y(alu_out_5_) );
NOR2X1 NOR2X1_1379 ( .A(_5160_), .B(_5159_), .Y(_3280_) );
INVX1 INVX1_1287 ( .A(_3280_), .Y(_3281_) );
INVX1 INVX1_1288 ( .A(_5183_), .Y(_3282_) );
OAI21X1 OAI21X1_3594 ( .A(_3234_), .B(_5170_), .C(_3282_), .Y(_3283_) );
INVX1 INVX1_1289 ( .A(_3283_), .Y(_3284_) );
OAI21X1 OAI21X1_3595 ( .A(_10734__5_), .B(_10728__5_), .C(_3258_), .Y(_3285_) );
OAI21X1 OAI21X1_3596 ( .A(_5179_), .B(_5862_), .C(_3285_), .Y(_3286_) );
MUX2X1 MUX2X1_281 ( .A(_3286_), .B(_3284_), .S(_3223__bF_buf1), .Y(_3287_) );
AND2X2 AND2X2_230 ( .A(_3287_), .B(_3281_), .Y(_3288_) );
OAI21X1 OAI21X1_3597 ( .A(_3287_), .B(_3281_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0), .Y(_3289_) );
OAI21X1 OAI21X1_3598 ( .A(_3161_), .B(_10728__2_bF_buf0_), .C(_3262_), .Y(_3290_) );
INVX1 INVX1_1290 ( .A(_3290_), .Y(_3291_) );
NAND2X1 NAND2X1_1149 ( .A(_10728__2_bF_buf4_), .B(_3163_), .Y(_3292_) );
OAI21X1 OAI21X1_3599 ( .A(_3169_), .B(_10728__2_bF_buf3_), .C(_3292_), .Y(_3293_) );
NAND2X1 NAND2X1_1150 ( .A(_5856__bF_buf1), .B(_3293_), .Y(_3294_) );
OAI21X1 OAI21X1_3600 ( .A(_5856__bF_buf0), .B(_3291_), .C(_3294_), .Y(_3295_) );
NAND2X1 NAND2X1_1151 ( .A(_5131__bF_buf2), .B(_3154_), .Y(_3296_) );
AOI21X1 AOI21X1_995 ( .A(_10728__2_bF_buf2_), .B(_3158_), .C(_10728__3_bF_buf1_), .Y(_3297_) );
NAND2X1 NAND2X1_1152 ( .A(_10728__2_bF_buf1_), .B(_3171_), .Y(_3298_) );
OAI21X1 OAI21X1_3601 ( .A(_10728__2_bF_buf0_), .B(_3157_), .C(_3298_), .Y(_3299_) );
AOI22X1 AOI22X1_160 ( .A(_3296_), .B(_3297_), .C(_3299_), .D(_10728__3_bF_buf0_), .Y(_3300_) );
AOI21X1 AOI21X1_996 ( .A(_5859__bF_buf3), .B(_3300_), .C(_3041_), .Y(_3301_) );
OAI21X1 OAI21X1_3602 ( .A(_5859__bF_buf2), .B(_3295_), .C(_3301_), .Y(_3302_) );
OAI22X1 OAI22X1_291 ( .A(_3007__bF_buf2), .B(_5158_), .C(_5160_), .D(_3005__bF_buf3), .Y(_3303_) );
AOI21X1 AOI21X1_997 ( .A(_3011__bF_buf4), .B(_3280_), .C(_3303_), .Y(_3304_) );
AND2X2 AND2X2_231 ( .A(_3302_), .B(_3304_), .Y(_3305_) );
OAI21X1 OAI21X1_3603 ( .A(_3288_), .B(_3289_), .C(_3305_), .Y(alu_out_6_) );
NOR2X1 NOR2X1_1380 ( .A(_3280_), .B(_3284_), .Y(_3306_) );
OAI21X1 OAI21X1_3604 ( .A(_3306_), .B(_5175_), .C(instr_sub_bF_buf4), .Y(_3307_) );
NAND2X1 NAND2X1_1153 ( .A(_3280_), .B(_3286_), .Y(_3308_) );
OAI21X1 OAI21X1_3605 ( .A(_5174_), .B(_5926_), .C(_3308_), .Y(_3309_) );
OAI21X1 OAI21X1_3606 ( .A(_3309_), .B(instr_sub_bF_buf3), .C(_3307_), .Y(_3310_) );
AND2X2 AND2X2_232 ( .A(_3310_), .B(_5157_), .Y(_3311_) );
OAI21X1 OAI21X1_3607 ( .A(_3310_), .B(_5157_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .Y(_3312_) );
OAI22X1 OAI22X1_292 ( .A(_3007__bF_buf1), .B(_5153_), .C(_5155_), .D(_3005__bF_buf2), .Y(_3313_) );
AOI21X1 AOI21X1_998 ( .A(_3011__bF_buf3), .B(_5156_), .C(_3313_), .Y(_3314_) );
NAND2X1 NAND2X1_1154 ( .A(_5131__bF_buf1), .B(_3199_), .Y(_3315_) );
OAI21X1 OAI21X1_3608 ( .A(_3191_), .B(_5131__bF_buf0), .C(_3315_), .Y(_3316_) );
NOR2X1 NOR2X1_1381 ( .A(_10728__2_bF_buf4_), .B(_3192_), .Y(_3317_) );
NAND2X1 NAND2X1_1155 ( .A(_10728__3_bF_buf4_), .B(_3079_), .Y(_3318_) );
OAI22X1 OAI22X1_293 ( .A(_3317_), .B(_3318_), .C(_3316_), .D(_10728__3_bF_buf3_), .Y(_3319_) );
INVX1 INVX1_1291 ( .A(_3319_), .Y(_3320_) );
NAND2X1 NAND2X1_1156 ( .A(_10728__2_bF_buf3_), .B(_3217_), .Y(_3321_) );
OAI21X1 OAI21X1_3609 ( .A(_3210_), .B(_10728__2_bF_buf2_), .C(_3321_), .Y(_3322_) );
NAND2X1 NAND2X1_1157 ( .A(_10728__2_bF_buf1_), .B(_3202_), .Y(_3323_) );
OAI21X1 OAI21X1_3610 ( .A(_3215_), .B(_10728__2_bF_buf0_), .C(_3323_), .Y(_3324_) );
MUX2X1 MUX2X1_282 ( .A(_3324_), .B(_3322_), .S(_10728__3_bF_buf2_), .Y(_3325_) );
AOI21X1 AOI21X1_999 ( .A(_5859__bF_buf1), .B(_3325_), .C(_3041_), .Y(_3326_) );
OAI21X1 OAI21X1_3611 ( .A(_5859__bF_buf0), .B(_3320_), .C(_3326_), .Y(_3327_) );
AND2X2 AND2X2_233 ( .A(_3327_), .B(_3314_), .Y(_3328_) );
OAI21X1 OAI21X1_3612 ( .A(_3311_), .B(_3312_), .C(_3328_), .Y(alu_out_7_) );
OAI21X1 OAI21X1_3613 ( .A(_5162_), .B(_5167_), .C(_5163_), .Y(_3329_) );
OAI21X1 OAI21X1_3614 ( .A(_5155_), .B(_5158_), .C(_5153_), .Y(_3330_) );
NOR2X1 NOR2X1_1382 ( .A(_5157_), .B(_3281_), .Y(_3331_) );
AOI21X1 AOI21X1_1000 ( .A(_3329_), .B(_3331_), .C(_3330_), .Y(_3332_) );
NOR2X1 NOR2X1_1383 ( .A(_5166_), .B(_3257_), .Y(_3333_) );
NAND3X1 NAND3X1_111 ( .A(_3333_), .B(_3331_), .C(_3237_), .Y(_3334_) );
NAND2X1 NAND2X1_1158 ( .A(_3332_), .B(_3334_), .Y(_3335_) );
INVX1 INVX1_1292 ( .A(_3335_), .Y(_3336_) );
NAND2X1 NAND2X1_1159 ( .A(_3223__bF_buf0), .B(_3336_), .Y(_3337_) );
OAI21X1 OAI21X1_3615 ( .A(_3223__bF_buf3), .B(_5185_), .C(_3337_), .Y(_3338_) );
AND2X2 AND2X2_234 ( .A(_3338_), .B(_5114_), .Y(_3339_) );
OAI21X1 OAI21X1_3616 ( .A(_3338_), .B(_5114_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3), .Y(_3340_) );
NOR2X1 NOR2X1_1384 ( .A(_10728__3_bF_buf1_), .B(_3024_), .Y(_3341_) );
OAI21X1 OAI21X1_3617 ( .A(_3072_), .B(_5856__bF_buf4), .C(_5859__bF_buf4), .Y(_3342_) );
NAND2X1 NAND2X1_1160 ( .A(_10728__3_bF_buf0_), .B(_3193_), .Y(_3343_) );
OAI21X1 OAI21X1_3618 ( .A(_3058_), .B(_10728__3_bF_buf4_), .C(_3343_), .Y(_3344_) );
NAND2X1 NAND2X1_1161 ( .A(_10728__4_bF_buf4_), .B(_3344_), .Y(_3345_) );
OAI21X1 OAI21X1_3619 ( .A(_3341_), .B(_3342_), .C(_3345_), .Y(_3346_) );
NOR2X1 NOR2X1_1385 ( .A(_3010_), .B(_5114_), .Y(_3347_) );
OAI22X1 OAI22X1_294 ( .A(_3007__bF_buf0), .B(_5110_), .C(_5112_), .D(_3005__bF_buf1), .Y(_3348_) );
OR2X2 OR2X2_46 ( .A(_3347_), .B(_3348_), .Y(_3349_) );
AOI21X1 AOI21X1_1001 ( .A(_3040_), .B(_3346_), .C(_3349_), .Y(_3350_) );
OAI21X1 OAI21X1_3620 ( .A(_3339_), .B(_3340_), .C(_3350_), .Y(alu_out_8_) );
NOR2X1 NOR2X1_1386 ( .A(_5106_), .B(_5109_), .Y(_3351_) );
INVX1 INVX1_1293 ( .A(_3351_), .Y(_3352_) );
NOR2X1 NOR2X1_1387 ( .A(_5114_), .B(_3336_), .Y(_3353_) );
OAI21X1 OAI21X1_3621 ( .A(_5187_), .B(_6051_), .C(_3223__bF_buf2), .Y(_3354_) );
NOR2X1 NOR2X1_1388 ( .A(_5113_), .B(_5185_), .Y(_3355_) );
OAI21X1 OAI21X1_3622 ( .A(_3355_), .B(_5188_), .C(instr_sub_bF_buf2), .Y(_3356_) );
OAI21X1 OAI21X1_3623 ( .A(_3353_), .B(_3354_), .C(_3356_), .Y(_3357_) );
AND2X2 AND2X2_235 ( .A(_3357_), .B(_3352_), .Y(_3358_) );
OAI21X1 OAI21X1_3624 ( .A(_3357_), .B(_3352_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2), .Y(_3359_) );
OAI21X1 OAI21X1_3625 ( .A(_3091_), .B(_10728__3_bF_buf3_), .C(_3343_), .Y(_3360_) );
NAND2X1 NAND2X1_1162 ( .A(_5856__bF_buf3), .B(_3127_), .Y(_3361_) );
OAI21X1 OAI21X1_3626 ( .A(_5856__bF_buf2), .B(_3107_), .C(_3361_), .Y(_3362_) );
AOI21X1 AOI21X1_1002 ( .A(_5859__bF_buf3), .B(_3362_), .C(_3041_), .Y(_3363_) );
OAI21X1 OAI21X1_3627 ( .A(_5859__bF_buf2), .B(_3360_), .C(_3363_), .Y(_3364_) );
INVX1 INVX1_1294 ( .A(_5109_), .Y(_3365_) );
OAI22X1 OAI22X1_295 ( .A(_5106_), .B(_3005__bF_buf0), .C(_3365_), .D(_3007__bF_buf4), .Y(_3366_) );
AOI21X1 AOI21X1_1003 ( .A(_3011__bF_buf2), .B(_3351_), .C(_3366_), .Y(_3367_) );
AND2X2 AND2X2_236 ( .A(_3364_), .B(_3367_), .Y(_3368_) );
OAI21X1 OAI21X1_3628 ( .A(_3358_), .B(_3359_), .C(_3368_), .Y(alu_out_9_) );
NOR2X1 NOR2X1_1389 ( .A(_5124_), .B(_5123_), .Y(_3369_) );
INVX1 INVX1_1295 ( .A(_3369_), .Y(_3370_) );
OR2X2 OR2X2_47 ( .A(_5185_), .B(_5115_), .Y(_3371_) );
AND2X2 AND2X2_237 ( .A(_3371_), .B(_5191_), .Y(_3372_) );
OAI21X1 OAI21X1_3629 ( .A(_5106_), .B(_5110_), .C(_3365_), .Y(_3373_) );
NOR2X1 NOR2X1_1390 ( .A(_5114_), .B(_3352_), .Y(_3374_) );
AOI21X1 AOI21X1_1004 ( .A(_3374_), .B(_3335_), .C(_3373_), .Y(_3375_) );
NOR2X1 NOR2X1_1391 ( .A(instr_sub_bF_buf1), .B(_3375_), .Y(_3376_) );
AOI21X1 AOI21X1_1005 ( .A(instr_sub_bF_buf0), .B(_3372_), .C(_3376_), .Y(_3377_) );
AND2X2 AND2X2_238 ( .A(_3377_), .B(_3370_), .Y(_3378_) );
OAI21X1 OAI21X1_3630 ( .A(_3377_), .B(_3370_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1), .Y(_3379_) );
MUX2X1 MUX2X1_283 ( .A(_3173_), .B(_3159_), .S(_10728__3_bF_buf2_), .Y(_3380_) );
OAI21X1 OAI21X1_3631 ( .A(_3166_), .B(_10728__3_bF_buf1_), .C(_3343_), .Y(_3381_) );
NAND2X1 NAND2X1_1163 ( .A(_10728__4_bF_buf3_), .B(_3381_), .Y(_3382_) );
OAI21X1 OAI21X1_3632 ( .A(_10728__4_bF_buf2_), .B(_3380_), .C(_3382_), .Y(_3383_) );
NOR2X1 NOR2X1_1392 ( .A(_3010_), .B(_3370_), .Y(_3384_) );
OAI21X1 OAI21X1_3633 ( .A(instr_andi), .B(instr_and), .C(_5123_), .Y(_3385_) );
OAI21X1 OAI21X1_3634 ( .A(_5124_), .B(_3005__bF_buf4), .C(_3385_), .Y(_3386_) );
OR2X2 OR2X2_48 ( .A(_3384_), .B(_3386_), .Y(_3387_) );
AOI21X1 AOI21X1_1006 ( .A(_3040_), .B(_3383_), .C(_3387_), .Y(_3388_) );
OAI21X1 OAI21X1_3635 ( .A(_3378_), .B(_3379_), .C(_3388_), .Y(alu_out_10_) );
NOR2X1 NOR2X1_1393 ( .A(_3369_), .B(_3372_), .Y(_3389_) );
AOI21X1 AOI21X1_1007 ( .A(_10734__10_), .B(_5122_), .C(_3389_), .Y(_3390_) );
NOR2X1 NOR2X1_1394 ( .A(instr_sub_bF_buf4), .B(_5123_), .Y(_3391_) );
OAI21X1 OAI21X1_3636 ( .A(_3375_), .B(_5124_), .C(_3391_), .Y(_3392_) );
OAI21X1 OAI21X1_3637 ( .A(_3390_), .B(_3223__bF_buf1), .C(_3392_), .Y(_3393_) );
AND2X2 AND2X2_239 ( .A(_3393_), .B(_5120_), .Y(_3394_) );
OAI21X1 OAI21X1_3638 ( .A(_3393_), .B(_5120_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0), .Y(_3395_) );
NOR2X1 NOR2X1_1395 ( .A(_5116_), .B(_3007__bF_buf3), .Y(_3396_) );
AOI21X1 AOI21X1_1008 ( .A(_5119_), .B(_3006_), .C(_3396_), .Y(_3397_) );
OAI21X1 OAI21X1_3639 ( .A(_5120_), .B(_3010_), .C(_3397_), .Y(_3398_) );
OAI21X1 OAI21X1_3640 ( .A(_3196_), .B(_10728__3_bF_buf0_), .C(_3343_), .Y(_3399_) );
NOR2X1 NOR2X1_1396 ( .A(_5859__bF_buf1), .B(_3399_), .Y(_3400_) );
INVX1 INVX1_1296 ( .A(_3204_), .Y(_3401_) );
NAND2X1 NAND2X1_1164 ( .A(_5856__bF_buf1), .B(_3219_), .Y(_3402_) );
OAI21X1 OAI21X1_3641 ( .A(_3401_), .B(_5856__bF_buf0), .C(_3402_), .Y(_3403_) );
OAI21X1 OAI21X1_3642 ( .A(_3403_), .B(_10728__4_bF_buf1_), .C(_3040_), .Y(_3404_) );
NOR2X1 NOR2X1_1397 ( .A(_3400_), .B(_3404_), .Y(_3405_) );
NOR2X1 NOR2X1_1398 ( .A(_3398_), .B(_3405_), .Y(_3406_) );
OAI21X1 OAI21X1_3643 ( .A(_3394_), .B(_3395_), .C(_3406_), .Y(alu_out_11_) );
NOR2X1 NOR2X1_1399 ( .A(_5120_), .B(_3370_), .Y(_3407_) );
NAND2X1 NAND2X1_1165 ( .A(_3374_), .B(_3407_), .Y(_3408_) );
INVX1 INVX1_1297 ( .A(_3408_), .Y(_3409_) );
NAND2X1 NAND2X1_1166 ( .A(_3373_), .B(_3407_), .Y(_3410_) );
INVX1 INVX1_1298 ( .A(_3410_), .Y(_3411_) );
INVX1 INVX1_1299 ( .A(_5123_), .Y(_3412_) );
OAI21X1 OAI21X1_3644 ( .A(_5120_), .B(_3412_), .C(_5116_), .Y(_3413_) );
OR2X2 OR2X2_49 ( .A(_3411_), .B(_3413_), .Y(_3414_) );
AOI21X1 AOI21X1_1009 ( .A(_3409_), .B(_3335_), .C(_3414_), .Y(_3415_) );
INVX1 INVX1_1300 ( .A(_3415_), .Y(_3416_) );
NAND2X1 NAND2X1_1167 ( .A(_3223__bF_buf0), .B(_3416_), .Y(_3417_) );
OAI21X1 OAI21X1_3645 ( .A(_5185_), .B(_5127_), .C(_5194_), .Y(_3418_) );
OAI21X1 OAI21X1_3646 ( .A(_3223__bF_buf3), .B(_3418_), .C(_3417_), .Y(_3419_) );
AOI21X1 AOI21X1_1010 ( .A(_5098_), .B(_3419_), .C(_3184_), .Y(_3420_) );
OAI21X1 OAI21X1_3647 ( .A(_5098_), .B(_3419_), .C(_3420_), .Y(_3421_) );
OAI22X1 OAI22X1_296 ( .A(_3007__bF_buf2), .B(_5095_), .C(_5097_), .D(_3005__bF_buf3), .Y(_3422_) );
AOI21X1 AOI21X1_1011 ( .A(_3011__bF_buf1), .B(_5098_), .C(_3422_), .Y(_3423_) );
OAI21X1 OAI21X1_3648 ( .A(_3246_), .B(_10728__3_bF_buf4_), .C(_3343_), .Y(_3424_) );
MUX2X1 MUX2X1_284 ( .A(_3247_), .B(_3243_), .S(_10728__3_bF_buf3_), .Y(_3425_) );
AOI21X1 AOI21X1_1012 ( .A(_5859__bF_buf0), .B(_3425_), .C(_3041_), .Y(_3426_) );
OAI21X1 OAI21X1_3649 ( .A(_5859__bF_buf4), .B(_3424_), .C(_3426_), .Y(_3427_) );
NAND3X1 NAND3X1_112 ( .A(_3423_), .B(_3427_), .C(_3421_), .Y(alu_out_12_) );
NOR2X1 NOR2X1_1400 ( .A(_5102_), .B(_5101_), .Y(_3428_) );
INVX1 INVX1_1301 ( .A(_3428_), .Y(_3429_) );
OAI21X1 OAI21X1_3650 ( .A(_5096_), .B(_5097_), .C(_3418_), .Y(_3430_) );
INVX1 INVX1_1302 ( .A(_3430_), .Y(_3431_) );
OAI21X1 OAI21X1_3651 ( .A(_3431_), .B(_5198_), .C(instr_sub_bF_buf3), .Y(_3432_) );
OAI21X1 OAI21X1_3652 ( .A(_3415_), .B(_5097_), .C(_5095_), .Y(_3433_) );
OAI21X1 OAI21X1_3653 ( .A(instr_sub_bF_buf2), .B(_3433_), .C(_3432_), .Y(_3434_) );
AND2X2 AND2X2_240 ( .A(_3434_), .B(_3429_), .Y(_3435_) );
OAI21X1 OAI21X1_3654 ( .A(_3434_), .B(_3429_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .Y(_3436_) );
OAI21X1 OAI21X1_3655 ( .A(_3264_), .B(_10728__3_bF_buf2_), .C(_3343_), .Y(_3437_) );
MUX2X1 MUX2X1_285 ( .A(_3267_), .B(_3271_), .S(_10728__3_bF_buf1_), .Y(_3438_) );
AOI21X1 AOI21X1_1013 ( .A(_5859__bF_buf3), .B(_3438_), .C(_3041_), .Y(_3439_) );
OAI21X1 OAI21X1_3656 ( .A(_5859__bF_buf2), .B(_3437_), .C(_3439_), .Y(_3440_) );
OAI22X1 OAI22X1_297 ( .A(_3007__bF_buf1), .B(_5100_), .C(_5102_), .D(_3005__bF_buf2), .Y(_3441_) );
AOI21X1 AOI21X1_1014 ( .A(_3011__bF_buf0), .B(_3428_), .C(_3441_), .Y(_3442_) );
AND2X2 AND2X2_241 ( .A(_3440_), .B(_3442_), .Y(_3443_) );
OAI21X1 OAI21X1_3657 ( .A(_3435_), .B(_3436_), .C(_3443_), .Y(alu_out_13_) );
NOR2X1 NOR2X1_1401 ( .A(_5093_), .B(_5092_), .Y(_3444_) );
INVX1 INVX1_1303 ( .A(_3444_), .Y(_3445_) );
OAI21X1 OAI21X1_3658 ( .A(_3430_), .B(_3428_), .C(_5201_), .Y(_3446_) );
NOR2X1 NOR2X1_1402 ( .A(_3223__bF_buf2), .B(_3446_), .Y(_3447_) );
NOR2X1 NOR2X1_1403 ( .A(_5099_), .B(_3429_), .Y(_3448_) );
OAI21X1 OAI21X1_3659 ( .A(_5102_), .B(_5095_), .C(_5100_), .Y(_3449_) );
AOI21X1 AOI21X1_1015 ( .A(_3448_), .B(_3416_), .C(_3449_), .Y(_3450_) );
NOR2X1 NOR2X1_1404 ( .A(instr_sub_bF_buf1), .B(_3450_), .Y(_3451_) );
NOR2X1 NOR2X1_1405 ( .A(_3451_), .B(_3447_), .Y(_3452_) );
AND2X2 AND2X2_242 ( .A(_3452_), .B(_3445_), .Y(_3453_) );
OAI21X1 OAI21X1_3660 ( .A(_3452_), .B(_3445_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3), .Y(_3454_) );
OAI21X1 OAI21X1_3661 ( .A(instr_andi), .B(instr_and), .C(_5092_), .Y(_3455_) );
NOR2X1 NOR2X1_1406 ( .A(_10728__3_bF_buf0_), .B(_3299_), .Y(_3456_) );
OAI21X1 OAI21X1_3662 ( .A(_3293_), .B(_5856__bF_buf4), .C(_5859__bF_buf1), .Y(_3457_) );
OAI21X1 OAI21X1_3663 ( .A(_3290_), .B(_10728__3_bF_buf4_), .C(_3318_), .Y(_3458_) );
OAI22X1 OAI22X1_298 ( .A(_3458_), .B(_5859__bF_buf0), .C(_3457_), .D(_3456_), .Y(_3459_) );
OAI22X1 OAI22X1_299 ( .A(_5093_), .B(_3005__bF_buf1), .C(_3445_), .D(_3010_), .Y(_3460_) );
AOI21X1 AOI21X1_1016 ( .A(_3040_), .B(_3459_), .C(_3460_), .Y(_3461_) );
AND2X2 AND2X2_243 ( .A(_3461_), .B(_3455_), .Y(_3462_) );
OAI21X1 OAI21X1_3664 ( .A(_3453_), .B(_3454_), .C(_3462_), .Y(alu_out_14_) );
AND2X2 AND2X2_244 ( .A(_3446_), .B(_3445_), .Y(_3463_) );
OAI21X1 OAI21X1_3665 ( .A(_3463_), .B(_5204_), .C(instr_sub_bF_buf0), .Y(_3464_) );
OAI21X1 OAI21X1_3666 ( .A(_3450_), .B(_3445_), .C(_5091_), .Y(_3465_) );
OAI21X1 OAI21X1_3667 ( .A(instr_sub_bF_buf4), .B(_3465_), .C(_3464_), .Y(_3466_) );
AND2X2 AND2X2_245 ( .A(_3466_), .B(_5090_), .Y(_3467_) );
OAI21X1 OAI21X1_3668 ( .A(_3466_), .B(_5090_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2), .Y(_3468_) );
MUX2X1 MUX2X1_286 ( .A(_3324_), .B(_3316_), .S(_5856__bF_buf3), .Y(_3469_) );
OAI21X1 OAI21X1_3669 ( .A(_3317_), .B(_3193_), .C(_5856__bF_buf2), .Y(_3470_) );
OAI21X1 OAI21X1_3670 ( .A(_5856__bF_buf1), .B(_3079_), .C(_3470_), .Y(_3471_) );
NAND2X1 NAND2X1_1168 ( .A(_10728__4_bF_buf0_), .B(_3471_), .Y(_3472_) );
OAI21X1 OAI21X1_3671 ( .A(_3469_), .B(_10728__4_bF_buf4_), .C(_3472_), .Y(_3473_) );
INVX1 INVX1_1304 ( .A(_5086_), .Y(_3474_) );
AOI22X1 AOI22X1_161 ( .A(_3006_), .B(_5089_), .C(_3474_), .D(_3008_), .Y(_3475_) );
OAI21X1 OAI21X1_3672 ( .A(_5090_), .B(_3010_), .C(_3475_), .Y(_3476_) );
AOI21X1 AOI21X1_1017 ( .A(_3040_), .B(_3473_), .C(_3476_), .Y(_3477_) );
OAI21X1 OAI21X1_3673 ( .A(_3467_), .B(_3468_), .C(_3477_), .Y(alu_out_15_) );
NOR2X1 NOR2X1_1407 ( .A(_5207_), .B(_5186_), .Y(_3478_) );
NAND2X1 NAND2X1_1169 ( .A(instr_sub_bF_buf3), .B(_3478_), .Y(_3479_) );
INVX1 INVX1_1305 ( .A(_3449_), .Y(_3480_) );
OR2X2 OR2X2_50 ( .A(_3445_), .B(_5090_), .Y(_3481_) );
AOI21X1 AOI21X1_1018 ( .A(_5089_), .B(_5092_), .C(_3474_), .Y(_3482_) );
OAI21X1 OAI21X1_3674 ( .A(_3481_), .B(_3480_), .C(_3482_), .Y(_3483_) );
INVX1 INVX1_1306 ( .A(_3448_), .Y(_3484_) );
NOR2X1 NOR2X1_1408 ( .A(_3481_), .B(_3484_), .Y(_3485_) );
AOI21X1 AOI21X1_1019 ( .A(_3485_), .B(_3414_), .C(_3483_), .Y(_3486_) );
NAND2X1 NAND2X1_1170 ( .A(_3485_), .B(_3409_), .Y(_3487_) );
OAI21X1 OAI21X1_3675 ( .A(_3336_), .B(_3487_), .C(_3486_), .Y(_3488_) );
INVX1 INVX1_1307 ( .A(_3488_), .Y(_3489_) );
OAI21X1 OAI21X1_3676 ( .A(instr_sub_bF_buf2), .B(_3489_), .C(_3479_), .Y(_3490_) );
AOI21X1 AOI21X1_1020 ( .A(_5055_), .B(_3490_), .C(_3184_), .Y(_3491_) );
OAI21X1 OAI21X1_3677 ( .A(_5055_), .B(_3490_), .C(_3491_), .Y(_3492_) );
INVX1 INVX1_1308 ( .A(_5053_), .Y(_3493_) );
OAI22X1 OAI22X1_300 ( .A(_5054_), .B(_3005__bF_buf0), .C(_3493_), .D(_3007__bF_buf0), .Y(_3494_) );
AOI21X1 AOI21X1_1021 ( .A(_3011__bF_buf4), .B(_5055_), .C(_3494_), .Y(_3495_) );
OAI21X1 OAI21X1_3678 ( .A(_5859__bF_buf4), .B(_3193_), .C(_3040_), .Y(_3496_) );
INVX1 INVX1_1309 ( .A(_3496_), .Y(_3497_) );
NAND2X1 NAND2X1_1171 ( .A(_5859__bF_buf3), .B(_3073_), .Y(_3498_) );
NAND2X1 NAND2X1_1172 ( .A(_3497_), .B(_3498_), .Y(_3499_) );
NAND3X1 NAND3X1_113 ( .A(_3495_), .B(_3499_), .C(_3492_), .Y(alu_out_16_) );
OAI21X1 OAI21X1_3679 ( .A(_5186_), .B(_5207_), .C(_5056_), .Y(_3500_) );
OAI21X1 OAI21X1_3680 ( .A(_3489_), .B(_5056_), .C(_3493_), .Y(_3501_) );
AOI21X1 AOI21X1_1022 ( .A(_10734__16_), .B(_5052_), .C(_3223__bF_buf1), .Y(_3502_) );
AOI22X1 AOI22X1_162 ( .A(_3500_), .B(_3502_), .C(_3501_), .D(_3223__bF_buf0), .Y(_3503_) );
AND2X2 AND2X2_246 ( .A(_3503_), .B(_5062_), .Y(_3504_) );
OAI21X1 OAI21X1_3681 ( .A(_3503_), .B(_5062_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1), .Y(_3505_) );
OAI21X1 OAI21X1_3682 ( .A(_3109_), .B(_10728__4_bF_buf3_), .C(_3497_), .Y(_3506_) );
INVX1 INVX1_1310 ( .A(_5059_), .Y(_3507_) );
OAI22X1 OAI22X1_301 ( .A(_5060_), .B(_3005__bF_buf4), .C(_3507_), .D(_3007__bF_buf4), .Y(_3508_) );
AOI21X1 AOI21X1_1023 ( .A(_3011__bF_buf3), .B(_5061_), .C(_3508_), .Y(_3509_) );
AND2X2 AND2X2_247 ( .A(_3506_), .B(_3509_), .Y(_3510_) );
OAI21X1 OAI21X1_3683 ( .A(_3504_), .B(_3505_), .C(_3510_), .Y(alu_out_17_) );
INVX1 INVX1_1311 ( .A(_5049_), .Y(_3511_) );
NOR2X1 NOR2X1_1409 ( .A(_5061_), .B(_3500_), .Y(_3512_) );
NOR2X1 NOR2X1_1410 ( .A(_5211_), .B(_3512_), .Y(_3513_) );
NOR2X1 NOR2X1_1411 ( .A(_5056_), .B(_5062_), .Y(_3514_) );
INVX1 INVX1_1312 ( .A(_3514_), .Y(_3515_) );
OAI21X1 OAI21X1_3684 ( .A(_3493_), .B(_5060_), .C(_3507_), .Y(_3516_) );
INVX1 INVX1_1313 ( .A(_3516_), .Y(_3517_) );
OAI21X1 OAI21X1_3685 ( .A(_3489_), .B(_3515_), .C(_3517_), .Y(_3518_) );
MUX2X1 MUX2X1_287 ( .A(_3513_), .B(_3518_), .S(instr_sub_bF_buf1), .Y(_3519_) );
AND2X2 AND2X2_248 ( .A(_3519_), .B(_3511_), .Y(_3520_) );
OAI21X1 OAI21X1_3686 ( .A(_3519_), .B(_3511_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0), .Y(_3521_) );
OAI21X1 OAI21X1_3687 ( .A(_3175_), .B(_10728__4_bF_buf2_), .C(_3497_), .Y(_3522_) );
INVX1 INVX1_1314 ( .A(_5047_), .Y(_3523_) );
OAI22X1 OAI22X1_302 ( .A(_5048_), .B(_3005__bF_buf3), .C(_3523_), .D(_3007__bF_buf3), .Y(_3524_) );
AOI21X1 AOI21X1_1024 ( .A(_3011__bF_buf2), .B(_5049_), .C(_3524_), .Y(_3525_) );
AND2X2 AND2X2_249 ( .A(_3522_), .B(_3525_), .Y(_3526_) );
OAI21X1 OAI21X1_3688 ( .A(_3520_), .B(_3521_), .C(_3526_), .Y(alu_out_18_) );
OAI21X1 OAI21X1_3689 ( .A(_3512_), .B(_5211_), .C(_3511_), .Y(_3527_) );
OAI21X1 OAI21X1_3690 ( .A(_5045_), .B(_10735__18_), .C(_3527_), .Y(_3528_) );
NAND2X1 NAND2X1_1173 ( .A(instr_sub_bF_buf0), .B(_3528_), .Y(_3529_) );
AOI21X1 AOI21X1_1025 ( .A(_5049_), .B(_3518_), .C(_5047_), .Y(_3530_) );
NAND2X1 NAND2X1_1174 ( .A(_3223__bF_buf3), .B(_3530_), .Y(_3531_) );
AOI21X1 AOI21X1_1026 ( .A(_3531_), .B(_3529_), .C(_5044_), .Y(_3532_) );
NAND2X1 NAND2X1_1175 ( .A(_3531_), .B(_3529_), .Y(_3533_) );
OAI21X1 OAI21X1_3691 ( .A(_3533_), .B(_5212_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .Y(_3534_) );
OAI21X1 OAI21X1_3692 ( .A(_3206_), .B(_10728__4_bF_buf1_), .C(_3497_), .Y(_3535_) );
INVX1 INVX1_1315 ( .A(_5042_), .Y(_3536_) );
OAI22X1 OAI22X1_303 ( .A(_5043_), .B(_3005__bF_buf2), .C(_3536_), .D(_3007__bF_buf2), .Y(_3537_) );
AOI21X1 AOI21X1_1027 ( .A(_3011__bF_buf1), .B(_5044_), .C(_3537_), .Y(_3538_) );
AND2X2 AND2X2_250 ( .A(_3535_), .B(_3538_), .Y(_3539_) );
OAI21X1 OAI21X1_3693 ( .A(_3534_), .B(_3532_), .C(_3539_), .Y(alu_out_19_) );
INVX1 INVX1_1316 ( .A(_5076_), .Y(_3540_) );
NOR2X1 NOR2X1_1412 ( .A(_5212_), .B(_3511_), .Y(_3541_) );
NAND2X1 NAND2X1_1176 ( .A(_3541_), .B(_3514_), .Y(_3542_) );
INVX1 INVX1_1317 ( .A(_3542_), .Y(_3543_) );
OAI21X1 OAI21X1_3694 ( .A(_3523_), .B(_5043_), .C(_3536_), .Y(_3544_) );
AOI21X1 AOI21X1_1028 ( .A(_3516_), .B(_3541_), .C(_3544_), .Y(_3545_) );
INVX1 INVX1_1318 ( .A(_3545_), .Y(_3546_) );
AOI21X1 AOI21X1_1029 ( .A(_3543_), .B(_3488_), .C(_3546_), .Y(_3547_) );
NOR2X1 NOR2X1_1413 ( .A(instr_sub_bF_buf4), .B(_3547_), .Y(_3548_) );
OAI21X1 OAI21X1_3695 ( .A(_3478_), .B(_5063_), .C(_5215_), .Y(_3549_) );
NOR2X1 NOR2X1_1414 ( .A(_3223__bF_buf2), .B(_3549_), .Y(_3550_) );
NOR2X1 NOR2X1_1415 ( .A(_3548_), .B(_3550_), .Y(_3551_) );
AND2X2 AND2X2_251 ( .A(_3551_), .B(_3540_), .Y(_3552_) );
OAI21X1 OAI21X1_3696 ( .A(_3551_), .B(_3540_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3), .Y(_3553_) );
OAI21X1 OAI21X1_3697 ( .A(_3249_), .B(_10728__4_bF_buf0_), .C(_3497_), .Y(_3554_) );
OAI22X1 OAI22X1_304 ( .A(_3007__bF_buf1), .B(_5073_), .C(_5075_), .D(_3005__bF_buf1), .Y(_3555_) );
AOI21X1 AOI21X1_1030 ( .A(_3011__bF_buf0), .B(_5076_), .C(_3555_), .Y(_3556_) );
AND2X2 AND2X2_252 ( .A(_3554_), .B(_3556_), .Y(_3557_) );
OAI21X1 OAI21X1_3698 ( .A(_3552_), .B(_3553_), .C(_3557_), .Y(alu_out_20_) );
INVX1 INVX1_1319 ( .A(_5080_), .Y(_3558_) );
OAI21X1 OAI21X1_3699 ( .A(_3547_), .B(_3540_), .C(_5073_), .Y(_3559_) );
AOI21X1 AOI21X1_1031 ( .A(_3540_), .B(_3549_), .C(_5219_), .Y(_3560_) );
MUX2X1 MUX2X1_288 ( .A(_3560_), .B(_3559_), .S(instr_sub_bF_buf3), .Y(_3561_) );
AND2X2 AND2X2_253 ( .A(_3561_), .B(_3558_), .Y(_3562_) );
OAI21X1 OAI21X1_3700 ( .A(_3561_), .B(_3558_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2), .Y(_3563_) );
OAI21X1 OAI21X1_3701 ( .A(_3269_), .B(_10728__4_bF_buf4_), .C(_3497_), .Y(_3564_) );
OAI22X1 OAI22X1_305 ( .A(_3007__bF_buf0), .B(_5077_), .C(_5079_), .D(_3005__bF_buf0), .Y(_3565_) );
AOI21X1 AOI21X1_1032 ( .A(_3011__bF_buf4), .B(_5080_), .C(_3565_), .Y(_3566_) );
AND2X2 AND2X2_254 ( .A(_3564_), .B(_3566_), .Y(_3567_) );
OAI21X1 OAI21X1_3702 ( .A(_3562_), .B(_3563_), .C(_3567_), .Y(alu_out_21_) );
AOI21X1 AOI21X1_1033 ( .A(_5081_), .B(_3549_), .C(_5221_), .Y(_3568_) );
NAND2X1 NAND2X1_1177 ( .A(instr_sub_bF_buf2), .B(_3568_), .Y(_3569_) );
NOR2X1 NOR2X1_1416 ( .A(_3540_), .B(_3558_), .Y(_3570_) );
INVX1 INVX1_1320 ( .A(_3570_), .Y(_3571_) );
OAI21X1 OAI21X1_3703 ( .A(_5079_), .B(_5073_), .C(_5077_), .Y(_3572_) );
INVX1 INVX1_1321 ( .A(_3572_), .Y(_3573_) );
OAI21X1 OAI21X1_3704 ( .A(_3547_), .B(_3571_), .C(_3573_), .Y(_3574_) );
NAND2X1 NAND2X1_1178 ( .A(_3223__bF_buf1), .B(_3574_), .Y(_3575_) );
NAND2X1 NAND2X1_1179 ( .A(_3575_), .B(_3569_), .Y(_3576_) );
XNOR2X1 XNOR2X1_58 ( .A(_3576_), .B(_5071_), .Y(_3577_) );
OAI21X1 OAI21X1_3705 ( .A(_3295_), .B(_10728__4_bF_buf3_), .C(_3497_), .Y(_3578_) );
OAI22X1 OAI22X1_306 ( .A(_3007__bF_buf4), .B(_5068_), .C(_5070_), .D(_3005__bF_buf4), .Y(_3579_) );
AOI21X1 AOI21X1_1034 ( .A(_3011__bF_buf3), .B(_5071_), .C(_3579_), .Y(_3580_) );
AND2X2 AND2X2_255 ( .A(_3578_), .B(_3580_), .Y(_3581_) );
OAI21X1 OAI21X1_3706 ( .A(_3577_), .B(_3184_), .C(_3581_), .Y(alu_out_22_) );
OAI21X1 OAI21X1_3707 ( .A(_3568_), .B(_5071_), .C(_5225_), .Y(_3582_) );
AOI21X1 AOI21X1_1035 ( .A(_5071_), .B(_3574_), .C(_5069_), .Y(_3583_) );
MUX2X1 MUX2X1_289 ( .A(_3582_), .B(_3583_), .S(instr_sub_bF_buf1), .Y(_3584_) );
AND2X2 AND2X2_256 ( .A(_3584_), .B(_5067_), .Y(_3585_) );
OAI21X1 OAI21X1_3708 ( .A(_3584_), .B(_5067_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1), .Y(_3586_) );
OAI21X1 OAI21X1_3709 ( .A(_3320_), .B(_10728__4_bF_buf2_), .C(_3497_), .Y(_3587_) );
OAI22X1 OAI22X1_307 ( .A(_3007__bF_buf3), .B(_5064_), .C(_5066_), .D(_3005__bF_buf3), .Y(_3588_) );
AOI21X1 AOI21X1_1036 ( .A(_3011__bF_buf2), .B(_5067_), .C(_3588_), .Y(_3589_) );
AND2X2 AND2X2_257 ( .A(_3587_), .B(_3589_), .Y(_3590_) );
OAI21X1 OAI21X1_3710 ( .A(_3585_), .B(_3586_), .C(_3590_), .Y(alu_out_23_) );
INVX1 INVX1_1322 ( .A(_5036_), .Y(_3591_) );
AND2X2 AND2X2_258 ( .A(_5067_), .B(_5071_), .Y(_3592_) );
OAI21X1 OAI21X1_3711 ( .A(_5066_), .B(_5068_), .C(_5064_), .Y(_3593_) );
AOI21X1 AOI21X1_1037 ( .A(_3572_), .B(_3592_), .C(_3593_), .Y(_3594_) );
NAND2X1 NAND2X1_1180 ( .A(_3592_), .B(_3570_), .Y(_3595_) );
OAI21X1 OAI21X1_3712 ( .A(_3545_), .B(_3595_), .C(_3594_), .Y(_3596_) );
NOR2X1 NOR2X1_1417 ( .A(_3595_), .B(_3542_), .Y(_3597_) );
AOI21X1 AOI21X1_1038 ( .A(_3597_), .B(_3488_), .C(_3596_), .Y(_3598_) );
INVX1 INVX1_1323 ( .A(_3598_), .Y(_3599_) );
INVX1 INVX1_1324 ( .A(_5229_), .Y(_3600_) );
OAI21X1 OAI21X1_3713 ( .A(_5186_), .B(_5207_), .C(_5083_), .Y(_3601_) );
AND2X2 AND2X2_259 ( .A(_3601_), .B(_3600_), .Y(_3602_) );
MUX2X1 MUX2X1_290 ( .A(_3599_), .B(_3602_), .S(_3223__bF_buf0), .Y(_3603_) );
AND2X2 AND2X2_260 ( .A(_3603_), .B(_3591_), .Y(_3604_) );
OAI21X1 OAI21X1_3714 ( .A(_3603_), .B(_3591_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0), .Y(_3605_) );
OAI21X1 OAI21X1_3715 ( .A(_3344_), .B(_10728__4_bF_buf1_), .C(_3497_), .Y(_3606_) );
INVX1 INVX1_1325 ( .A(_5034_), .Y(_3607_) );
OAI22X1 OAI22X1_308 ( .A(_5035_), .B(_3005__bF_buf2), .C(_3607_), .D(_3007__bF_buf2), .Y(_3608_) );
AOI21X1 AOI21X1_1039 ( .A(_3011__bF_buf1), .B(_5036_), .C(_3608_), .Y(_3609_) );
AND2X2 AND2X2_261 ( .A(_3606_), .B(_3609_), .Y(_3610_) );
OAI21X1 OAI21X1_3716 ( .A(_3604_), .B(_3605_), .C(_3610_), .Y(alu_out_24_) );
INVX1 INVX1_1326 ( .A(_5031_), .Y(_3611_) );
OAI21X1 OAI21X1_3717 ( .A(_3598_), .B(_5035_), .C(_3607_), .Y(_3612_) );
NOR2X1 NOR2X1_1418 ( .A(_5036_), .B(_3602_), .Y(_3613_) );
NOR2X1 NOR2X1_1419 ( .A(_5230_), .B(_3613_), .Y(_3614_) );
MUX2X1 MUX2X1_291 ( .A(_3614_), .B(_3612_), .S(instr_sub_bF_buf0), .Y(_3615_) );
AND2X2 AND2X2_262 ( .A(_3615_), .B(_3611_), .Y(_3616_) );
OAI21X1 OAI21X1_3718 ( .A(_3615_), .B(_3611_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .Y(_3617_) );
OAI21X1 OAI21X1_3719 ( .A(_3360_), .B(_10728__4_bF_buf0_), .C(_3497_), .Y(_3618_) );
INVX1 INVX1_1327 ( .A(_5030_), .Y(_3619_) );
AOI22X1 AOI22X1_163 ( .A(_3619_), .B(_3006_), .C(_5031_), .D(_3011__bF_buf0), .Y(_3620_) );
NAND2X1 NAND2X1_1181 ( .A(_3620_), .B(_3618_), .Y(_3621_) );
AOI21X1 AOI21X1_1040 ( .A(_5029_), .B(_3008_), .C(_3621_), .Y(_3622_) );
OAI21X1 OAI21X1_3720 ( .A(_3616_), .B(_3617_), .C(_3622_), .Y(alu_out_25_) );
INVX1 INVX1_1328 ( .A(_5037_), .Y(_3623_) );
INVX1 INVX1_1329 ( .A(_5232_), .Y(_3624_) );
OAI21X1 OAI21X1_3721 ( .A(_3602_), .B(_3623_), .C(_3624_), .Y(_3625_) );
NOR2X1 NOR2X1_1420 ( .A(_3611_), .B(_3591_), .Y(_3626_) );
INVX1 INVX1_1330 ( .A(_3626_), .Y(_3627_) );
AOI21X1 AOI21X1_1041 ( .A(_3619_), .B(_5034_), .C(_5029_), .Y(_3628_) );
OAI21X1 OAI21X1_3722 ( .A(_3598_), .B(_3627_), .C(_3628_), .Y(_3629_) );
NAND2X1 NAND2X1_1182 ( .A(_3223__bF_buf3), .B(_3629_), .Y(_3630_) );
OAI21X1 OAI21X1_3723 ( .A(_3625_), .B(_3223__bF_buf2), .C(_3630_), .Y(_3631_) );
AOI21X1 AOI21X1_1042 ( .A(_5025_), .B(_3631_), .C(_3184_), .Y(_3632_) );
OAI21X1 OAI21X1_3724 ( .A(_5025_), .B(_3631_), .C(_3632_), .Y(_3633_) );
OAI21X1 OAI21X1_3725 ( .A(_3381_), .B(_10728__4_bF_buf4_), .C(_3497_), .Y(_3634_) );
INVX1 INVX1_1331 ( .A(_5023_), .Y(_3635_) );
OAI22X1 OAI22X1_309 ( .A(_5024_), .B(_3005__bF_buf1), .C(_3635_), .D(_3007__bF_buf1), .Y(_3636_) );
AOI21X1 AOI21X1_1043 ( .A(_3011__bF_buf4), .B(_5025_), .C(_3636_), .Y(_3637_) );
NAND3X1 NAND3X1_114 ( .A(_3634_), .B(_3637_), .C(_3633_), .Y(alu_out_26_) );
INVX1 INVX1_1332 ( .A(_5020_), .Y(_3638_) );
INVX1 INVX1_1333 ( .A(_5025_), .Y(_3639_) );
AOI21X1 AOI21X1_1044 ( .A(_3639_), .B(_3625_), .C(_5235_), .Y(_3640_) );
OAI21X1 OAI21X1_3726 ( .A(_10734__26_), .B(_10735__26_), .C(_3629_), .Y(_3641_) );
OAI21X1 OAI21X1_3727 ( .A(_5021_), .B(_5022_), .C(_3641_), .Y(_3642_) );
MUX2X1 MUX2X1_292 ( .A(_3642_), .B(_3640_), .S(_3223__bF_buf1), .Y(_3643_) );
AND2X2 AND2X2_263 ( .A(_3643_), .B(_3638_), .Y(_3644_) );
OAI21X1 OAI21X1_3728 ( .A(_3643_), .B(_3638_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf3), .Y(_3645_) );
OAI21X1 OAI21X1_3729 ( .A(_3399_), .B(_10728__4_bF_buf3_), .C(_3497_), .Y(_3646_) );
INVX1 INVX1_1334 ( .A(_5018_), .Y(_3647_) );
OAI22X1 OAI22X1_310 ( .A(_5019_), .B(_3005__bF_buf0), .C(_3647_), .D(_3007__bF_buf0), .Y(_3648_) );
AOI21X1 AOI21X1_1045 ( .A(_3011__bF_buf3), .B(_5020_), .C(_3648_), .Y(_3649_) );
AND2X2 AND2X2_264 ( .A(_3646_), .B(_3649_), .Y(_3650_) );
OAI21X1 OAI21X1_3730 ( .A(_3644_), .B(_3645_), .C(_3650_), .Y(alu_out_27_) );
INVX1 INVX1_1335 ( .A(_5008_), .Y(_3651_) );
NOR2X1 NOR2X1_1421 ( .A(_3638_), .B(_3639_), .Y(_3652_) );
INVX1 INVX1_1336 ( .A(_3652_), .Y(_3653_) );
NOR2X1 NOR2X1_1422 ( .A(_3627_), .B(_3653_), .Y(_3654_) );
INVX1 INVX1_1337 ( .A(_3654_), .Y(_3655_) );
OAI21X1 OAI21X1_3731 ( .A(_3635_), .B(_5019_), .C(_3647_), .Y(_3656_) );
INVX1 INVX1_1338 ( .A(_3656_), .Y(_3657_) );
OAI21X1 OAI21X1_3732 ( .A(_3653_), .B(_3628_), .C(_3657_), .Y(_3658_) );
INVX1 INVX1_1339 ( .A(_3658_), .Y(_3659_) );
OAI21X1 OAI21X1_3733 ( .A(_3598_), .B(_3655_), .C(_3659_), .Y(_3660_) );
OAI21X1 OAI21X1_3734 ( .A(_3602_), .B(_5038_), .C(_5239_), .Y(_3661_) );
NOR2X1 NOR2X1_1423 ( .A(_3223__bF_buf0), .B(_3661_), .Y(_3662_) );
AOI21X1 AOI21X1_1046 ( .A(_3223__bF_buf3), .B(_3660_), .C(_3662_), .Y(_3663_) );
AND2X2 AND2X2_265 ( .A(_3663_), .B(_3651_), .Y(_3664_) );
OAI21X1 OAI21X1_3735 ( .A(_3663_), .B(_3651_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf2), .Y(_3665_) );
OAI21X1 OAI21X1_3736 ( .A(_3424_), .B(_10728__4_bF_buf2_), .C(_3497_), .Y(_3666_) );
INVX1 INVX1_1340 ( .A(_5006_), .Y(_3667_) );
OAI22X1 OAI22X1_311 ( .A(_5007_), .B(_3005__bF_buf4), .C(_3667_), .D(_3007__bF_buf4), .Y(_3668_) );
AOI21X1 AOI21X1_1047 ( .A(_3011__bF_buf2), .B(_5008_), .C(_3668_), .Y(_3669_) );
AND2X2 AND2X2_266 ( .A(_3666_), .B(_3669_), .Y(_3670_) );
OAI21X1 OAI21X1_3737 ( .A(_3664_), .B(_3665_), .C(_3670_), .Y(alu_out_28_) );
INVX1 INVX1_1341 ( .A(_5013_), .Y(_3671_) );
INVX1 INVX1_1342 ( .A(_3660_), .Y(_3672_) );
OAI21X1 OAI21X1_3738 ( .A(_3672_), .B(_5007_), .C(_3667_), .Y(_3673_) );
AOI21X1 AOI21X1_1048 ( .A(_3651_), .B(_3661_), .C(_5240_), .Y(_3674_) );
MUX2X1 MUX2X1_293 ( .A(_3673_), .B(_3674_), .S(_3223__bF_buf2), .Y(_3675_) );
AND2X2 AND2X2_267 ( .A(_3675_), .B(_3671_), .Y(_3676_) );
OAI21X1 OAI21X1_3739 ( .A(_3675_), .B(_3671_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf1), .Y(_3677_) );
OR2X2 OR2X2_51 ( .A(_3437_), .B(_10728__4_bF_buf1_), .Y(_3678_) );
AOI22X1 AOI22X1_164 ( .A(_5011_), .B(_3008_), .C(_5013_), .D(_3011__bF_buf1), .Y(_3679_) );
OAI21X1 OAI21X1_3740 ( .A(_5012_), .B(_3005__bF_buf3), .C(_3679_), .Y(_3680_) );
AOI21X1 AOI21X1_1049 ( .A(_3497_), .B(_3678_), .C(_3680_), .Y(_3681_) );
OAI21X1 OAI21X1_3741 ( .A(_3676_), .B(_3677_), .C(_3681_), .Y(alu_out_29_) );
INVX1 INVX1_1343 ( .A(_5002_), .Y(_3682_) );
INVX1 INVX1_1344 ( .A(_5242_), .Y(_3683_) );
AOI21X1 AOI21X1_1050 ( .A(_3600_), .B(_3601_), .C(_5038_), .Y(_3684_) );
OAI21X1 OAI21X1_3742 ( .A(_3684_), .B(_5238_), .C(_5014_), .Y(_3685_) );
AND2X2 AND2X2_268 ( .A(_3685_), .B(_3683_), .Y(_3686_) );
NOR2X1 NOR2X1_1424 ( .A(_3651_), .B(_3671_), .Y(_3687_) );
AOI21X1 AOI21X1_1051 ( .A(_5006_), .B(_5013_), .C(_5011_), .Y(_3688_) );
INVX1 INVX1_1345 ( .A(_3688_), .Y(_3689_) );
AOI21X1 AOI21X1_1052 ( .A(_3687_), .B(_3660_), .C(_3689_), .Y(_3690_) );
NOR2X1 NOR2X1_1425 ( .A(instr_sub_bF_buf4), .B(_3690_), .Y(_3691_) );
AOI21X1 AOI21X1_1053 ( .A(instr_sub_bF_buf3), .B(_3686_), .C(_3691_), .Y(_3692_) );
AND2X2 AND2X2_269 ( .A(_3692_), .B(_3682_), .Y(_3693_) );
OAI21X1 OAI21X1_3743 ( .A(_3692_), .B(_3682_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf0), .Y(_3694_) );
NAND2X1 NAND2X1_1183 ( .A(_5859__bF_buf2), .B(_3458_), .Y(_3695_) );
INVX1 INVX1_1346 ( .A(_5001_), .Y(_3696_) );
AOI22X1 AOI22X1_165 ( .A(_3696_), .B(_3006_), .C(_5000_), .D(_3008_), .Y(_3697_) );
OAI21X1 OAI21X1_3744 ( .A(_3682_), .B(_3010_), .C(_3697_), .Y(_3698_) );
AOI21X1 AOI21X1_1054 ( .A(_3497_), .B(_3695_), .C(_3698_), .Y(_3699_) );
OAI21X1 OAI21X1_3745 ( .A(_3693_), .B(_3694_), .C(_3699_), .Y(alu_out_30_) );
NOR2X1 NOR2X1_1426 ( .A(instr_sub_bF_buf2), .B(_5000_), .Y(_3700_) );
OAI21X1 OAI21X1_3746 ( .A(_3690_), .B(_5001_), .C(_3700_), .Y(_3701_) );
AOI21X1 AOI21X1_1055 ( .A(_3683_), .B(_3685_), .C(_5002_), .Y(_3702_) );
OAI21X1 OAI21X1_3747 ( .A(_3702_), .B(_5243_), .C(instr_sub_bF_buf1), .Y(_3703_) );
AOI21X1 AOI21X1_1056 ( .A(_3701_), .B(_3703_), .C(_4996_), .Y(_3704_) );
NAND2X1 NAND2X1_1184 ( .A(_3701_), .B(_3703_), .Y(_3705_) );
OAI21X1 OAI21X1_3748 ( .A(_3705_), .B(_4997_), .C(is_lui_auipc_jal_jalr_addi_add_sub_bF_buf4), .Y(_3706_) );
AOI22X1 AOI22X1_166 ( .A(_4995_), .B(_3008_), .C(_4996_), .D(_3011__bF_buf0), .Y(_3707_) );
OAI21X1 OAI21X1_3749 ( .A(_4993_), .B(_3005__bF_buf2), .C(_3707_), .Y(_3708_) );
AOI21X1 AOI21X1_1057 ( .A(_3471_), .B(_3497_), .C(_3708_), .Y(_3709_) );
OAI21X1 OAI21X1_3750 ( .A(_3706_), .B(_3704_), .C(_3709_), .Y(alu_out_31_) );
INVX1 INVX1_1347 ( .A(_4668_), .Y(_3710_) );
NAND2X1 NAND2X1_1185 ( .A(_5270_), .B(_3710_), .Y(_3711_) );
NAND2X1 NAND2X1_1186 ( .A(cpuregs_10_[0]), .B(_3711__bF_buf7), .Y(_3712_) );
OAI21X1 OAI21X1_3751 ( .A(_4925__bF_buf1), .B(_3711__bF_buf6), .C(_3712_), .Y(_731_) );
NAND2X1 NAND2X1_1187 ( .A(cpuregs_10_[1]), .B(_3711__bF_buf5), .Y(_3713_) );
OAI21X1 OAI21X1_3752 ( .A(_4933__bF_buf1), .B(_3711__bF_buf4), .C(_3713_), .Y(_732_) );
NAND2X1 NAND2X1_1188 ( .A(cpuregs_10_[2]), .B(_3711__bF_buf3), .Y(_3714_) );
OAI21X1 OAI21X1_3753 ( .A(_4940__bF_buf1), .B(_3711__bF_buf2), .C(_3714_), .Y(_733_) );
NAND2X1 NAND2X1_1189 ( .A(cpuregs_10_[3]), .B(_3711__bF_buf1), .Y(_3715_) );
OAI21X1 OAI21X1_3754 ( .A(_4948__bF_buf1), .B(_3711__bF_buf0), .C(_3715_), .Y(_734_) );
NAND2X1 NAND2X1_1190 ( .A(cpuregs_10_[4]), .B(_3711__bF_buf7), .Y(_3716_) );
OAI21X1 OAI21X1_3755 ( .A(_4955__bF_buf2), .B(_3711__bF_buf6), .C(_3716_), .Y(_735_) );
NAND2X1 NAND2X1_1191 ( .A(cpuregs_10_[5]), .B(_3711__bF_buf5), .Y(_3717_) );
OAI21X1 OAI21X1_3756 ( .A(_4654__bF_buf1), .B(_3711__bF_buf4), .C(_3717_), .Y(_736_) );
NAND2X1 NAND2X1_1192 ( .A(cpuregs_10_[6]), .B(_3711__bF_buf3), .Y(_3718_) );
OAI21X1 OAI21X1_3757 ( .A(_4664__bF_buf1), .B(_3711__bF_buf2), .C(_3718_), .Y(_737_) );
NAND2X1 NAND2X1_1193 ( .A(cpuregs_10_[7]), .B(_3711__bF_buf1), .Y(_3719_) );
OAI21X1 OAI21X1_3758 ( .A(_4677__bF_buf0), .B(_3711__bF_buf0), .C(_3719_), .Y(_738_) );
NAND2X1 NAND2X1_1194 ( .A(cpuregs_10_[8]), .B(_3711__bF_buf7), .Y(_3720_) );
OAI21X1 OAI21X1_3759 ( .A(_4685__bF_buf1), .B(_3711__bF_buf6), .C(_3720_), .Y(_739_) );
NAND2X1 NAND2X1_1195 ( .A(cpuregs_10_[9]), .B(_3711__bF_buf5), .Y(_3721_) );
OAI21X1 OAI21X1_3760 ( .A(_4696__bF_buf0), .B(_3711__bF_buf4), .C(_3721_), .Y(_740_) );
NAND2X1 NAND2X1_1196 ( .A(cpuregs_10_[10]), .B(_3711__bF_buf3), .Y(_3722_) );
OAI21X1 OAI21X1_3761 ( .A(_4703__bF_buf0), .B(_3711__bF_buf2), .C(_3722_), .Y(_741_) );
NAND2X1 NAND2X1_1197 ( .A(cpuregs_10_[11]), .B(_3711__bF_buf1), .Y(_3723_) );
OAI21X1 OAI21X1_3762 ( .A(_4713__bF_buf0), .B(_3711__bF_buf0), .C(_3723_), .Y(_742_) );
NAND2X1 NAND2X1_1198 ( .A(cpuregs_10_[12]), .B(_3711__bF_buf7), .Y(_3724_) );
OAI21X1 OAI21X1_3763 ( .A(_4722__bF_buf0), .B(_3711__bF_buf6), .C(_3724_), .Y(_743_) );
NAND2X1 NAND2X1_1199 ( .A(cpuregs_10_[13]), .B(_3711__bF_buf5), .Y(_3725_) );
OAI21X1 OAI21X1_3764 ( .A(_4731__bF_buf0), .B(_3711__bF_buf4), .C(_3725_), .Y(_744_) );
NAND2X1 NAND2X1_1200 ( .A(cpuregs_10_[14]), .B(_3711__bF_buf3), .Y(_3726_) );
OAI21X1 OAI21X1_3765 ( .A(_4740__bF_buf0), .B(_3711__bF_buf2), .C(_3726_), .Y(_745_) );
NAND2X1 NAND2X1_1201 ( .A(cpuregs_10_[15]), .B(_3711__bF_buf1), .Y(_3727_) );
OAI21X1 OAI21X1_3766 ( .A(_4747__bF_buf0), .B(_3711__bF_buf0), .C(_3727_), .Y(_746_) );
NAND2X1 NAND2X1_1202 ( .A(cpuregs_10_[16]), .B(_3711__bF_buf7), .Y(_3728_) );
OAI21X1 OAI21X1_3767 ( .A(_4755__bF_buf0), .B(_3711__bF_buf6), .C(_3728_), .Y(_747_) );
NAND2X1 NAND2X1_1203 ( .A(cpuregs_10_[17]), .B(_3711__bF_buf5), .Y(_3729_) );
OAI21X1 OAI21X1_3768 ( .A(_4763__bF_buf0), .B(_3711__bF_buf4), .C(_3729_), .Y(_748_) );
NAND2X1 NAND2X1_1204 ( .A(cpuregs_10_[18]), .B(_3711__bF_buf3), .Y(_3730_) );
OAI21X1 OAI21X1_3769 ( .A(_4783__bF_buf0), .B(_3711__bF_buf2), .C(_3730_), .Y(_749_) );
NAND2X1 NAND2X1_1205 ( .A(cpuregs_10_[19]), .B(_3711__bF_buf1), .Y(_3731_) );
OAI21X1 OAI21X1_3770 ( .A(_4793__bF_buf0), .B(_3711__bF_buf0), .C(_3731_), .Y(_750_) );
NAND2X1 NAND2X1_1206 ( .A(cpuregs_10_[20]), .B(_3711__bF_buf7), .Y(_3732_) );
OAI21X1 OAI21X1_3771 ( .A(_4806__bF_buf0), .B(_3711__bF_buf6), .C(_3732_), .Y(_751_) );
NAND2X1 NAND2X1_1207 ( .A(cpuregs_10_[21]), .B(_3711__bF_buf5), .Y(_3733_) );
OAI21X1 OAI21X1_3772 ( .A(_4816__bF_buf0), .B(_3711__bF_buf4), .C(_3733_), .Y(_752_) );
NAND2X1 NAND2X1_1208 ( .A(cpuregs_10_[22]), .B(_3711__bF_buf3), .Y(_3734_) );
OAI21X1 OAI21X1_3773 ( .A(_4824__bF_buf0), .B(_3711__bF_buf2), .C(_3734_), .Y(_753_) );
NAND2X1 NAND2X1_1209 ( .A(cpuregs_10_[23]), .B(_3711__bF_buf1), .Y(_3735_) );
OAI21X1 OAI21X1_3774 ( .A(_4833__bF_buf0), .B(_3711__bF_buf0), .C(_3735_), .Y(_754_) );
NAND2X1 NAND2X1_1210 ( .A(cpuregs_10_[24]), .B(_3711__bF_buf7), .Y(_3736_) );
OAI21X1 OAI21X1_3775 ( .A(_4845__bF_buf0), .B(_3711__bF_buf6), .C(_3736_), .Y(_755_) );
NAND2X1 NAND2X1_1211 ( .A(cpuregs_10_[25]), .B(_3711__bF_buf5), .Y(_3737_) );
OAI21X1 OAI21X1_3776 ( .A(_4854__bF_buf0), .B(_3711__bF_buf4), .C(_3737_), .Y(_756_) );
NAND2X1 NAND2X1_1212 ( .A(cpuregs_10_[26]), .B(_3711__bF_buf3), .Y(_3738_) );
OAI21X1 OAI21X1_3777 ( .A(_4863__bF_buf0), .B(_3711__bF_buf2), .C(_3738_), .Y(_757_) );
NAND2X1 NAND2X1_1213 ( .A(cpuregs_10_[27]), .B(_3711__bF_buf1), .Y(_3739_) );
OAI21X1 OAI21X1_3778 ( .A(_4871__bF_buf0), .B(_3711__bF_buf0), .C(_3739_), .Y(_758_) );
NAND2X1 NAND2X1_1214 ( .A(cpuregs_10_[28]), .B(_3711__bF_buf7), .Y(_3740_) );
OAI21X1 OAI21X1_3779 ( .A(_4884__bF_buf0), .B(_3711__bF_buf6), .C(_3740_), .Y(_759_) );
NAND2X1 NAND2X1_1215 ( .A(cpuregs_10_[29]), .B(_3711__bF_buf5), .Y(_3741_) );
OAI21X1 OAI21X1_3780 ( .A(_4893__bF_buf0), .B(_3711__bF_buf4), .C(_3741_), .Y(_760_) );
NAND2X1 NAND2X1_1216 ( .A(cpuregs_10_[30]), .B(_3711__bF_buf3), .Y(_3742_) );
OAI21X1 OAI21X1_3781 ( .A(_4901__bF_buf0), .B(_3711__bF_buf2), .C(_3742_), .Y(_761_) );
NAND2X1 NAND2X1_1217 ( .A(cpuregs_10_[31]), .B(_3711__bF_buf1), .Y(_3743_) );
OAI21X1 OAI21X1_3782 ( .A(_4910__bF_buf0), .B(_3711__bF_buf0), .C(_3743_), .Y(_762_) );
NOR2X1 NOR2X1_1427 ( .A(_5312_), .B(_4668_), .Y(_3744_) );
NOR2X1 NOR2X1_1428 ( .A(cpuregs_9_[0]), .B(_3744_), .Y(_3745_) );
AOI21X1 AOI21X1_1058 ( .A(_4925__bF_buf0), .B(_3744_), .C(_3745_), .Y(_763_) );
NAND2X1 NAND2X1_1218 ( .A(_5311_), .B(_4636_), .Y(_3746_) );
NOR2X1 NOR2X1_1429 ( .A(_3746__bF_buf3), .B(_4632__bF_buf6), .Y(_3747_) );
MUX2X1 MUX2X1_294 ( .A(_4933__bF_buf0), .B(_7669_), .S(_3747_), .Y(_764_) );
NOR2X1 NOR2X1_1430 ( .A(cpuregs_9_[2]), .B(_3744_), .Y(_3748_) );
AOI21X1 AOI21X1_1059 ( .A(_4940__bF_buf0), .B(_3744_), .C(_3748_), .Y(_765_) );
NOR2X1 NOR2X1_1431 ( .A(cpuregs_9_[3]), .B(_3744_), .Y(_3749_) );
AOI21X1 AOI21X1_1060 ( .A(_4948__bF_buf0), .B(_3744_), .C(_3749_), .Y(_766_) );
NOR2X1 NOR2X1_1432 ( .A(cpuregs_9_[4]), .B(_3744_), .Y(_3750_) );
AOI21X1 AOI21X1_1061 ( .A(_4955__bF_buf1), .B(_3744_), .C(_3750_), .Y(_767_) );
NAND2X1 NAND2X1_1219 ( .A(_3747_), .B(_4655_), .Y(_3751_) );
OAI21X1 OAI21X1_3783 ( .A(_5875_), .B(_3747_), .C(_3751_), .Y(_768_) );
NAND2X1 NAND2X1_1220 ( .A(_3747_), .B(_4665_), .Y(_3752_) );
OAI21X1 OAI21X1_3784 ( .A(_5939_), .B(_3747_), .C(_3752_), .Y(_769_) );
NAND2X1 NAND2X1_1221 ( .A(_3747_), .B(_2319_), .Y(_3753_) );
OAI21X1 OAI21X1_3785 ( .A(_5991_), .B(_3747_), .C(_3753_), .Y(_770_) );
NAND2X1 NAND2X1_1222 ( .A(_3747_), .B(_4686_), .Y(_3754_) );
OAI21X1 OAI21X1_3786 ( .A(_6070_), .B(_3747_), .C(_3754_), .Y(_771_) );
MUX2X1 MUX2X1_295 ( .A(_4696__bF_buf4), .B(_6127_), .S(_3744_), .Y(_772_) );
MUX2X1 MUX2X1_296 ( .A(_4703__bF_buf4), .B(_6177_), .S(_3744_), .Y(_773_) );
MUX2X1 MUX2X1_297 ( .A(_4713__bF_buf4), .B(_6256_), .S(_3744_), .Y(_774_) );
INVX1 INVX1_1348 ( .A(_3744_), .Y(_3755_) );
OAI21X1 OAI21X1_3787 ( .A(_4632__bF_buf5), .B(_3746__bF_buf2), .C(cpuregs_9_[12]), .Y(_3756_) );
OAI21X1 OAI21X1_3788 ( .A(_4722__bF_buf4), .B(_3755__bF_buf3), .C(_3756_), .Y(_775_) );
OAI21X1 OAI21X1_3789 ( .A(_4632__bF_buf4), .B(_3746__bF_buf1), .C(cpuregs_9_[13]), .Y(_3757_) );
OAI21X1 OAI21X1_3790 ( .A(_4731__bF_buf4), .B(_3755__bF_buf2), .C(_3757_), .Y(_776_) );
OAI21X1 OAI21X1_3791 ( .A(_4632__bF_buf3), .B(_3746__bF_buf0), .C(cpuregs_9_[14]), .Y(_3758_) );
OAI21X1 OAI21X1_3792 ( .A(_4740__bF_buf4), .B(_3755__bF_buf1), .C(_3758_), .Y(_777_) );
OAI21X1 OAI21X1_3793 ( .A(_4632__bF_buf2), .B(_3746__bF_buf3), .C(cpuregs_9_[15]), .Y(_3759_) );
OAI21X1 OAI21X1_3794 ( .A(_4747__bF_buf4), .B(_3755__bF_buf0), .C(_3759_), .Y(_778_) );
OAI21X1 OAI21X1_3795 ( .A(_4632__bF_buf1), .B(_3746__bF_buf2), .C(cpuregs_9_[16]), .Y(_3760_) );
OAI21X1 OAI21X1_3796 ( .A(_4755__bF_buf4), .B(_3755__bF_buf3), .C(_3760_), .Y(_779_) );
OAI21X1 OAI21X1_3797 ( .A(_4632__bF_buf0), .B(_3746__bF_buf1), .C(cpuregs_9_[17]), .Y(_3761_) );
OAI21X1 OAI21X1_3798 ( .A(_4763__bF_buf4), .B(_3755__bF_buf2), .C(_3761_), .Y(_780_) );
OAI21X1 OAI21X1_3799 ( .A(_4632__bF_buf8), .B(_3746__bF_buf0), .C(cpuregs_9_[18]), .Y(_3762_) );
OAI21X1 OAI21X1_3800 ( .A(_4783__bF_buf4), .B(_3755__bF_buf1), .C(_3762_), .Y(_781_) );
OAI21X1 OAI21X1_3801 ( .A(_4632__bF_buf7), .B(_3746__bF_buf3), .C(cpuregs_9_[19]), .Y(_3763_) );
OAI21X1 OAI21X1_3802 ( .A(_4793__bF_buf4), .B(_3755__bF_buf0), .C(_3763_), .Y(_782_) );
OAI21X1 OAI21X1_3803 ( .A(_4632__bF_buf6), .B(_3746__bF_buf2), .C(cpuregs_9_[20]), .Y(_3764_) );
OAI21X1 OAI21X1_3804 ( .A(_4806__bF_buf4), .B(_3755__bF_buf3), .C(_3764_), .Y(_783_) );
OAI21X1 OAI21X1_3805 ( .A(_4632__bF_buf5), .B(_3746__bF_buf1), .C(cpuregs_9_[21]), .Y(_3765_) );
OAI21X1 OAI21X1_3806 ( .A(_4816__bF_buf4), .B(_3755__bF_buf2), .C(_3765_), .Y(_784_) );
OAI21X1 OAI21X1_3807 ( .A(_4632__bF_buf4), .B(_3746__bF_buf0), .C(cpuregs_9_[22]), .Y(_3766_) );
OAI21X1 OAI21X1_3808 ( .A(_4824__bF_buf4), .B(_3755__bF_buf1), .C(_3766_), .Y(_785_) );
OAI21X1 OAI21X1_3809 ( .A(_4632__bF_buf3), .B(_3746__bF_buf3), .C(cpuregs_9_[23]), .Y(_3767_) );
OAI21X1 OAI21X1_3810 ( .A(_4833__bF_buf4), .B(_3755__bF_buf0), .C(_3767_), .Y(_786_) );
OAI21X1 OAI21X1_3811 ( .A(_4632__bF_buf2), .B(_3746__bF_buf2), .C(cpuregs_9_[24]), .Y(_3768_) );
OAI21X1 OAI21X1_3812 ( .A(_4845__bF_buf4), .B(_3755__bF_buf3), .C(_3768_), .Y(_787_) );
OAI21X1 OAI21X1_3813 ( .A(_4632__bF_buf1), .B(_3746__bF_buf1), .C(cpuregs_9_[25]), .Y(_3769_) );
OAI21X1 OAI21X1_3814 ( .A(_4854__bF_buf4), .B(_3755__bF_buf2), .C(_3769_), .Y(_788_) );
OAI21X1 OAI21X1_3815 ( .A(_4632__bF_buf0), .B(_3746__bF_buf0), .C(cpuregs_9_[26]), .Y(_3770_) );
OAI21X1 OAI21X1_3816 ( .A(_4863__bF_buf4), .B(_3755__bF_buf1), .C(_3770_), .Y(_789_) );
OAI21X1 OAI21X1_3817 ( .A(_4632__bF_buf8), .B(_3746__bF_buf3), .C(cpuregs_9_[27]), .Y(_3771_) );
OAI21X1 OAI21X1_3818 ( .A(_4871__bF_buf4), .B(_3755__bF_buf0), .C(_3771_), .Y(_790_) );
OAI21X1 OAI21X1_3819 ( .A(_4632__bF_buf7), .B(_3746__bF_buf2), .C(cpuregs_9_[28]), .Y(_3772_) );
OAI21X1 OAI21X1_3820 ( .A(_4884__bF_buf4), .B(_3755__bF_buf3), .C(_3772_), .Y(_791_) );
OAI21X1 OAI21X1_3821 ( .A(_4632__bF_buf6), .B(_3746__bF_buf1), .C(cpuregs_9_[29]), .Y(_3773_) );
OAI21X1 OAI21X1_3822 ( .A(_4893__bF_buf4), .B(_3755__bF_buf2), .C(_3773_), .Y(_792_) );
OAI21X1 OAI21X1_3823 ( .A(_4632__bF_buf5), .B(_3746__bF_buf0), .C(cpuregs_9_[30]), .Y(_3774_) );
OAI21X1 OAI21X1_3824 ( .A(_4901__bF_buf4), .B(_3755__bF_buf1), .C(_3774_), .Y(_793_) );
OAI21X1 OAI21X1_3825 ( .A(_4632__bF_buf4), .B(_3746__bF_buf3), .C(cpuregs_9_[31]), .Y(_3775_) );
OAI21X1 OAI21X1_3826 ( .A(_4910__bF_buf4), .B(_3755__bF_buf0), .C(_3775_), .Y(_794_) );
NAND2X1 NAND2X1_1223 ( .A(_4916_), .B(_3710_), .Y(_3776_) );
NAND2X1 NAND2X1_1224 ( .A(cpuregs_11_[0]), .B(_3776__bF_buf7), .Y(_3777_) );
OAI21X1 OAI21X1_3827 ( .A(_4925__bF_buf4), .B(_3776__bF_buf6), .C(_3777_), .Y(_795_) );
NAND2X1 NAND2X1_1225 ( .A(cpuregs_11_[1]), .B(_3776__bF_buf5), .Y(_3778_) );
OAI21X1 OAI21X1_3828 ( .A(_4933__bF_buf4), .B(_3776__bF_buf4), .C(_3778_), .Y(_796_) );
NAND2X1 NAND2X1_1226 ( .A(cpuregs_11_[2]), .B(_3776__bF_buf3), .Y(_3779_) );
OAI21X1 OAI21X1_3829 ( .A(_4940__bF_buf4), .B(_3776__bF_buf2), .C(_3779_), .Y(_797_) );
NAND2X1 NAND2X1_1227 ( .A(cpuregs_11_[3]), .B(_3776__bF_buf1), .Y(_3780_) );
OAI21X1 OAI21X1_3830 ( .A(_4948__bF_buf4), .B(_3776__bF_buf0), .C(_3780_), .Y(_798_) );
NAND2X1 NAND2X1_1228 ( .A(cpuregs_11_[4]), .B(_3776__bF_buf7), .Y(_3781_) );
OAI21X1 OAI21X1_3831 ( .A(_4955__bF_buf0), .B(_3776__bF_buf6), .C(_3781_), .Y(_799_) );
NAND2X1 NAND2X1_1229 ( .A(cpuregs_11_[5]), .B(_3776__bF_buf5), .Y(_3782_) );
OAI21X1 OAI21X1_3832 ( .A(_4654__bF_buf0), .B(_3776__bF_buf4), .C(_3782_), .Y(_800_) );
NAND2X1 NAND2X1_1230 ( .A(cpuregs_11_[6]), .B(_3776__bF_buf3), .Y(_3783_) );
OAI21X1 OAI21X1_3833 ( .A(_4664__bF_buf0), .B(_3776__bF_buf2), .C(_3783_), .Y(_801_) );
NAND2X1 NAND2X1_1231 ( .A(cpuregs_11_[7]), .B(_3776__bF_buf1), .Y(_3784_) );
OAI21X1 OAI21X1_3834 ( .A(_4677__bF_buf4), .B(_3776__bF_buf0), .C(_3784_), .Y(_802_) );
NAND2X1 NAND2X1_1232 ( .A(cpuregs_11_[8]), .B(_3776__bF_buf7), .Y(_3785_) );
OAI21X1 OAI21X1_3835 ( .A(_4685__bF_buf0), .B(_3776__bF_buf6), .C(_3785_), .Y(_803_) );
NAND2X1 NAND2X1_1233 ( .A(cpuregs_11_[9]), .B(_3776__bF_buf5), .Y(_3786_) );
OAI21X1 OAI21X1_3836 ( .A(_4696__bF_buf3), .B(_3776__bF_buf4), .C(_3786_), .Y(_804_) );
NAND2X1 NAND2X1_1234 ( .A(cpuregs_11_[10]), .B(_3776__bF_buf3), .Y(_3787_) );
OAI21X1 OAI21X1_3837 ( .A(_4703__bF_buf3), .B(_3776__bF_buf2), .C(_3787_), .Y(_805_) );
NAND2X1 NAND2X1_1235 ( .A(cpuregs_11_[11]), .B(_3776__bF_buf1), .Y(_3788_) );
OAI21X1 OAI21X1_3838 ( .A(_4713__bF_buf3), .B(_3776__bF_buf0), .C(_3788_), .Y(_806_) );
NAND2X1 NAND2X1_1236 ( .A(cpuregs_11_[12]), .B(_3776__bF_buf7), .Y(_3789_) );
OAI21X1 OAI21X1_3839 ( .A(_4722__bF_buf3), .B(_3776__bF_buf6), .C(_3789_), .Y(_807_) );
NAND2X1 NAND2X1_1237 ( .A(cpuregs_11_[13]), .B(_3776__bF_buf5), .Y(_3790_) );
OAI21X1 OAI21X1_3840 ( .A(_4731__bF_buf3), .B(_3776__bF_buf4), .C(_3790_), .Y(_808_) );
NAND2X1 NAND2X1_1238 ( .A(cpuregs_11_[14]), .B(_3776__bF_buf3), .Y(_3791_) );
OAI21X1 OAI21X1_3841 ( .A(_4740__bF_buf3), .B(_3776__bF_buf2), .C(_3791_), .Y(_809_) );
NAND2X1 NAND2X1_1239 ( .A(cpuregs_11_[15]), .B(_3776__bF_buf1), .Y(_3792_) );
OAI21X1 OAI21X1_3842 ( .A(_4747__bF_buf3), .B(_3776__bF_buf0), .C(_3792_), .Y(_810_) );
NAND2X1 NAND2X1_1240 ( .A(cpuregs_11_[16]), .B(_3776__bF_buf7), .Y(_3793_) );
OAI21X1 OAI21X1_3843 ( .A(_4755__bF_buf3), .B(_3776__bF_buf6), .C(_3793_), .Y(_811_) );
NAND2X1 NAND2X1_1241 ( .A(cpuregs_11_[17]), .B(_3776__bF_buf5), .Y(_3794_) );
OAI21X1 OAI21X1_3844 ( .A(_4763__bF_buf3), .B(_3776__bF_buf4), .C(_3794_), .Y(_812_) );
NAND2X1 NAND2X1_1242 ( .A(cpuregs_11_[18]), .B(_3776__bF_buf3), .Y(_3795_) );
OAI21X1 OAI21X1_3845 ( .A(_4783__bF_buf3), .B(_3776__bF_buf2), .C(_3795_), .Y(_813_) );
NAND2X1 NAND2X1_1243 ( .A(cpuregs_11_[19]), .B(_3776__bF_buf1), .Y(_3796_) );
OAI21X1 OAI21X1_3846 ( .A(_4793__bF_buf3), .B(_3776__bF_buf0), .C(_3796_), .Y(_814_) );
NAND2X1 NAND2X1_1244 ( .A(cpuregs_11_[20]), .B(_3776__bF_buf7), .Y(_3797_) );
OAI21X1 OAI21X1_3847 ( .A(_4806__bF_buf3), .B(_3776__bF_buf6), .C(_3797_), .Y(_815_) );
NAND2X1 NAND2X1_1245 ( .A(cpuregs_11_[21]), .B(_3776__bF_buf5), .Y(_3798_) );
OAI21X1 OAI21X1_3848 ( .A(_4816__bF_buf3), .B(_3776__bF_buf4), .C(_3798_), .Y(_816_) );
NAND2X1 NAND2X1_1246 ( .A(cpuregs_11_[22]), .B(_3776__bF_buf3), .Y(_3799_) );
OAI21X1 OAI21X1_3849 ( .A(_4824__bF_buf3), .B(_3776__bF_buf2), .C(_3799_), .Y(_817_) );
NAND2X1 NAND2X1_1247 ( .A(cpuregs_11_[23]), .B(_3776__bF_buf1), .Y(_3800_) );
OAI21X1 OAI21X1_3850 ( .A(_4833__bF_buf3), .B(_3776__bF_buf0), .C(_3800_), .Y(_818_) );
NAND2X1 NAND2X1_1248 ( .A(cpuregs_11_[24]), .B(_3776__bF_buf7), .Y(_3801_) );
OAI21X1 OAI21X1_3851 ( .A(_4845__bF_buf3), .B(_3776__bF_buf6), .C(_3801_), .Y(_819_) );
NAND2X1 NAND2X1_1249 ( .A(cpuregs_11_[25]), .B(_3776__bF_buf5), .Y(_3802_) );
OAI21X1 OAI21X1_3852 ( .A(_4854__bF_buf3), .B(_3776__bF_buf4), .C(_3802_), .Y(_820_) );
NAND2X1 NAND2X1_1250 ( .A(cpuregs_11_[26]), .B(_3776__bF_buf3), .Y(_3803_) );
OAI21X1 OAI21X1_3853 ( .A(_4863__bF_buf3), .B(_3776__bF_buf2), .C(_3803_), .Y(_821_) );
NAND2X1 NAND2X1_1251 ( .A(cpuregs_11_[27]), .B(_3776__bF_buf1), .Y(_3804_) );
OAI21X1 OAI21X1_3854 ( .A(_4871__bF_buf3), .B(_3776__bF_buf0), .C(_3804_), .Y(_822_) );
NAND2X1 NAND2X1_1252 ( .A(cpuregs_11_[28]), .B(_3776__bF_buf7), .Y(_3805_) );
OAI21X1 OAI21X1_3855 ( .A(_4884__bF_buf3), .B(_3776__bF_buf6), .C(_3805_), .Y(_823_) );
NAND2X1 NAND2X1_1253 ( .A(cpuregs_11_[29]), .B(_3776__bF_buf5), .Y(_3806_) );
OAI21X1 OAI21X1_3856 ( .A(_4893__bF_buf3), .B(_3776__bF_buf4), .C(_3806_), .Y(_824_) );
NAND2X1 NAND2X1_1254 ( .A(cpuregs_11_[30]), .B(_3776__bF_buf3), .Y(_3807_) );
OAI21X1 OAI21X1_3857 ( .A(_4901__bF_buf3), .B(_3776__bF_buf2), .C(_3807_), .Y(_825_) );
NAND2X1 NAND2X1_1255 ( .A(cpuregs_11_[31]), .B(_3776__bF_buf1), .Y(_3808_) );
OAI21X1 OAI21X1_3858 ( .A(_4910__bF_buf3), .B(_3776__bF_buf0), .C(_3808_), .Y(_826_) );
NOR2X1 NOR2X1_1433 ( .A(_2310__bF_buf5), .B(_5706__bF_buf8), .Y(_3809_) );
INVX1 INVX1_1349 ( .A(_3809_), .Y(_3810_) );
OAI21X1 OAI21X1_3859 ( .A(_5706__bF_buf7), .B(_2310__bF_buf4), .C(cpuregs_20_[0]), .Y(_3811_) );
OAI21X1 OAI21X1_3860 ( .A(_3810__bF_buf4), .B(_4925__bF_buf3), .C(_3811_), .Y(_827_) );
OAI21X1 OAI21X1_3861 ( .A(_5706__bF_buf6), .B(_2310__bF_buf3), .C(cpuregs_20_[1]), .Y(_3812_) );
OAI21X1 OAI21X1_3862 ( .A(_3810__bF_buf3), .B(_4933__bF_buf3), .C(_3812_), .Y(_828_) );
OAI21X1 OAI21X1_3863 ( .A(_5706__bF_buf5), .B(_2310__bF_buf2), .C(cpuregs_20_[2]), .Y(_3813_) );
OAI21X1 OAI21X1_3864 ( .A(_3810__bF_buf2), .B(_4940__bF_buf3), .C(_3813_), .Y(_829_) );
OAI21X1 OAI21X1_3865 ( .A(_5706__bF_buf4), .B(_2310__bF_buf1), .C(cpuregs_20_[3]), .Y(_3814_) );
OAI21X1 OAI21X1_3866 ( .A(_3810__bF_buf1), .B(_4948__bF_buf3), .C(_3814_), .Y(_830_) );
OAI21X1 OAI21X1_3867 ( .A(_5706__bF_buf3), .B(_2310__bF_buf0), .C(cpuregs_20_[4]), .Y(_3815_) );
OAI21X1 OAI21X1_3868 ( .A(_3810__bF_buf0), .B(_4955__bF_buf4), .C(_3815_), .Y(_831_) );
OAI21X1 OAI21X1_3869 ( .A(_5706__bF_buf2), .B(_2310__bF_buf7), .C(cpuregs_20_[5]), .Y(_3816_) );
OAI21X1 OAI21X1_3870 ( .A(_3810__bF_buf4), .B(_4654__bF_buf4), .C(_3816_), .Y(_832_) );
OAI21X1 OAI21X1_3871 ( .A(_5706__bF_buf1), .B(_2310__bF_buf6), .C(cpuregs_20_[6]), .Y(_3817_) );
OAI21X1 OAI21X1_3872 ( .A(_3810__bF_buf3), .B(_4664__bF_buf4), .C(_3817_), .Y(_833_) );
OAI21X1 OAI21X1_3873 ( .A(_5706__bF_buf0), .B(_2310__bF_buf5), .C(cpuregs_20_[7]), .Y(_3818_) );
OAI21X1 OAI21X1_3874 ( .A(_3810__bF_buf2), .B(_4677__bF_buf3), .C(_3818_), .Y(_834_) );
OAI21X1 OAI21X1_3875 ( .A(_5706__bF_buf11), .B(_2310__bF_buf4), .C(cpuregs_20_[8]), .Y(_3819_) );
OAI21X1 OAI21X1_3876 ( .A(_4685__bF_buf4), .B(_3810__bF_buf1), .C(_3819_), .Y(_835_) );
OAI21X1 OAI21X1_3877 ( .A(_5706__bF_buf10), .B(_2310__bF_buf3), .C(cpuregs_20_[9]), .Y(_3820_) );
OAI21X1 OAI21X1_3878 ( .A(_4696__bF_buf2), .B(_3810__bF_buf0), .C(_3820_), .Y(_836_) );
OAI21X1 OAI21X1_3879 ( .A(_5706__bF_buf9), .B(_2310__bF_buf2), .C(cpuregs_20_[10]), .Y(_3821_) );
OAI21X1 OAI21X1_3880 ( .A(_4703__bF_buf2), .B(_3810__bF_buf4), .C(_3821_), .Y(_837_) );
OAI21X1 OAI21X1_3881 ( .A(_5706__bF_buf8), .B(_2310__bF_buf1), .C(cpuregs_20_[11]), .Y(_3822_) );
OAI21X1 OAI21X1_3882 ( .A(_4713__bF_buf2), .B(_3810__bF_buf3), .C(_3822_), .Y(_838_) );
OAI21X1 OAI21X1_3883 ( .A(_5706__bF_buf7), .B(_2310__bF_buf0), .C(cpuregs_20_[12]), .Y(_3823_) );
OAI21X1 OAI21X1_3884 ( .A(_4722__bF_buf2), .B(_3810__bF_buf2), .C(_3823_), .Y(_839_) );
OAI21X1 OAI21X1_3885 ( .A(_5706__bF_buf6), .B(_2310__bF_buf7), .C(cpuregs_20_[13]), .Y(_3824_) );
OAI21X1 OAI21X1_3886 ( .A(_4731__bF_buf2), .B(_3810__bF_buf1), .C(_3824_), .Y(_840_) );
OAI21X1 OAI21X1_3887 ( .A(_5706__bF_buf5), .B(_2310__bF_buf6), .C(cpuregs_20_[14]), .Y(_3825_) );
OAI21X1 OAI21X1_3888 ( .A(_4740__bF_buf2), .B(_3810__bF_buf0), .C(_3825_), .Y(_841_) );
OAI21X1 OAI21X1_3889 ( .A(_5706__bF_buf4), .B(_2310__bF_buf5), .C(cpuregs_20_[15]), .Y(_3826_) );
OAI21X1 OAI21X1_3890 ( .A(_4747__bF_buf2), .B(_3810__bF_buf4), .C(_3826_), .Y(_842_) );
OAI21X1 OAI21X1_3891 ( .A(_5706__bF_buf3), .B(_2310__bF_buf4), .C(cpuregs_20_[16]), .Y(_3827_) );
OAI21X1 OAI21X1_3892 ( .A(_4755__bF_buf2), .B(_3810__bF_buf3), .C(_3827_), .Y(_843_) );
OAI21X1 OAI21X1_3893 ( .A(_5706__bF_buf2), .B(_2310__bF_buf3), .C(cpuregs_20_[17]), .Y(_3828_) );
OAI21X1 OAI21X1_3894 ( .A(_4763__bF_buf2), .B(_3810__bF_buf2), .C(_3828_), .Y(_844_) );
OAI21X1 OAI21X1_3895 ( .A(_5706__bF_buf1), .B(_2310__bF_buf2), .C(cpuregs_20_[18]), .Y(_3829_) );
OAI21X1 OAI21X1_3896 ( .A(_4783__bF_buf2), .B(_3810__bF_buf1), .C(_3829_), .Y(_845_) );
OAI21X1 OAI21X1_3897 ( .A(_5706__bF_buf0), .B(_2310__bF_buf1), .C(cpuregs_20_[19]), .Y(_3830_) );
OAI21X1 OAI21X1_3898 ( .A(_4793__bF_buf2), .B(_3810__bF_buf0), .C(_3830_), .Y(_846_) );
OAI21X1 OAI21X1_3899 ( .A(_5706__bF_buf11), .B(_2310__bF_buf0), .C(cpuregs_20_[20]), .Y(_3831_) );
OAI21X1 OAI21X1_3900 ( .A(_4806__bF_buf2), .B(_3810__bF_buf4), .C(_3831_), .Y(_847_) );
OAI21X1 OAI21X1_3901 ( .A(_5706__bF_buf10), .B(_2310__bF_buf7), .C(cpuregs_20_[21]), .Y(_3832_) );
OAI21X1 OAI21X1_3902 ( .A(_4816__bF_buf2), .B(_3810__bF_buf3), .C(_3832_), .Y(_848_) );
OAI21X1 OAI21X1_3903 ( .A(_5706__bF_buf9), .B(_2310__bF_buf6), .C(cpuregs_20_[22]), .Y(_3833_) );
OAI21X1 OAI21X1_3904 ( .A(_4824__bF_buf2), .B(_3810__bF_buf2), .C(_3833_), .Y(_849_) );
OAI21X1 OAI21X1_3905 ( .A(_5706__bF_buf8), .B(_2310__bF_buf5), .C(cpuregs_20_[23]), .Y(_3834_) );
OAI21X1 OAI21X1_3906 ( .A(_4833__bF_buf2), .B(_3810__bF_buf1), .C(_3834_), .Y(_850_) );
OAI21X1 OAI21X1_3907 ( .A(_5706__bF_buf7), .B(_2310__bF_buf4), .C(cpuregs_20_[24]), .Y(_3835_) );
OAI21X1 OAI21X1_3908 ( .A(_4845__bF_buf2), .B(_3810__bF_buf0), .C(_3835_), .Y(_851_) );
OAI21X1 OAI21X1_3909 ( .A(_5706__bF_buf6), .B(_2310__bF_buf3), .C(cpuregs_20_[25]), .Y(_3836_) );
OAI21X1 OAI21X1_3910 ( .A(_4854__bF_buf2), .B(_3810__bF_buf4), .C(_3836_), .Y(_852_) );
OAI21X1 OAI21X1_3911 ( .A(_5706__bF_buf5), .B(_2310__bF_buf2), .C(cpuregs_20_[26]), .Y(_3837_) );
OAI21X1 OAI21X1_3912 ( .A(_4863__bF_buf2), .B(_3810__bF_buf3), .C(_3837_), .Y(_853_) );
OAI21X1 OAI21X1_3913 ( .A(_5706__bF_buf4), .B(_2310__bF_buf1), .C(cpuregs_20_[27]), .Y(_3838_) );
OAI21X1 OAI21X1_3914 ( .A(_4871__bF_buf2), .B(_3810__bF_buf2), .C(_3838_), .Y(_854_) );
OAI21X1 OAI21X1_3915 ( .A(_5706__bF_buf3), .B(_2310__bF_buf0), .C(cpuregs_20_[28]), .Y(_3839_) );
OAI21X1 OAI21X1_3916 ( .A(_4884__bF_buf2), .B(_3810__bF_buf1), .C(_3839_), .Y(_855_) );
OAI21X1 OAI21X1_3917 ( .A(_5706__bF_buf2), .B(_2310__bF_buf7), .C(cpuregs_20_[29]), .Y(_3840_) );
OAI21X1 OAI21X1_3918 ( .A(_4893__bF_buf2), .B(_3810__bF_buf0), .C(_3840_), .Y(_856_) );
OAI21X1 OAI21X1_3919 ( .A(_5706__bF_buf1), .B(_2310__bF_buf6), .C(cpuregs_20_[30]), .Y(_3841_) );
OAI21X1 OAI21X1_3920 ( .A(_4901__bF_buf2), .B(_3810__bF_buf4), .C(_3841_), .Y(_857_) );
OAI21X1 OAI21X1_3921 ( .A(_5706__bF_buf0), .B(_2310__bF_buf5), .C(cpuregs_20_[31]), .Y(_3842_) );
OAI21X1 OAI21X1_3922 ( .A(_4910__bF_buf2), .B(_3810__bF_buf3), .C(_3842_), .Y(_858_) );
NOR2X1 NOR2X1_1434 ( .A(latched_rd_2_), .B(_2308_), .Y(_3843_) );
INVX1 INVX1_1350 ( .A(_3843_), .Y(_3844_) );
NOR2X1 NOR2X1_1435 ( .A(_3844__bF_buf8), .B(_4917__bF_buf9), .Y(_3845_) );
INVX1 INVX1_1351 ( .A(_3845_), .Y(_3846_) );
OAI21X1 OAI21X1_3923 ( .A(_4917__bF_buf8), .B(_3844__bF_buf7), .C(cpuregs_19_[0]), .Y(_3847_) );
OAI21X1 OAI21X1_3924 ( .A(_3846__bF_buf4), .B(_4925__bF_buf2), .C(_3847_), .Y(_859_) );
OAI21X1 OAI21X1_3925 ( .A(_4917__bF_buf7), .B(_3844__bF_buf6), .C(cpuregs_19_[1]), .Y(_3848_) );
OAI21X1 OAI21X1_3926 ( .A(_3846__bF_buf3), .B(_4933__bF_buf2), .C(_3848_), .Y(_860_) );
OAI21X1 OAI21X1_3927 ( .A(_4917__bF_buf6), .B(_3844__bF_buf5), .C(cpuregs_19_[2]), .Y(_3849_) );
OAI21X1 OAI21X1_3928 ( .A(_3846__bF_buf2), .B(_4940__bF_buf2), .C(_3849_), .Y(_861_) );
OAI21X1 OAI21X1_3929 ( .A(_4917__bF_buf5), .B(_3844__bF_buf4), .C(cpuregs_19_[3]), .Y(_3850_) );
OAI21X1 OAI21X1_3930 ( .A(_3846__bF_buf1), .B(_4948__bF_buf2), .C(_3850_), .Y(_862_) );
OAI21X1 OAI21X1_3931 ( .A(_4917__bF_buf4), .B(_3844__bF_buf3), .C(cpuregs_19_[4]), .Y(_3851_) );
OAI21X1 OAI21X1_3932 ( .A(_3846__bF_buf0), .B(_4955__bF_buf3), .C(_3851_), .Y(_863_) );
OAI21X1 OAI21X1_3933 ( .A(_4917__bF_buf3), .B(_3844__bF_buf2), .C(cpuregs_19_[5]), .Y(_3852_) );
OAI21X1 OAI21X1_3934 ( .A(_3846__bF_buf4), .B(_4654__bF_buf3), .C(_3852_), .Y(_864_) );
OAI21X1 OAI21X1_3935 ( .A(_4917__bF_buf2), .B(_3844__bF_buf1), .C(cpuregs_19_[6]), .Y(_3853_) );
OAI21X1 OAI21X1_3936 ( .A(_4664__bF_buf3), .B(_3846__bF_buf3), .C(_3853_), .Y(_865_) );
OAI21X1 OAI21X1_3937 ( .A(_4917__bF_buf1), .B(_3844__bF_buf0), .C(cpuregs_19_[7]), .Y(_3854_) );
OAI21X1 OAI21X1_3938 ( .A(_4677__bF_buf2), .B(_3846__bF_buf2), .C(_3854_), .Y(_866_) );
OAI21X1 OAI21X1_3939 ( .A(_4917__bF_buf0), .B(_3844__bF_buf8), .C(cpuregs_19_[8]), .Y(_3855_) );
OAI21X1 OAI21X1_3940 ( .A(_4685__bF_buf3), .B(_3846__bF_buf1), .C(_3855_), .Y(_867_) );
OAI21X1 OAI21X1_3941 ( .A(_4917__bF_buf10), .B(_3844__bF_buf7), .C(cpuregs_19_[9]), .Y(_3856_) );
OAI21X1 OAI21X1_3942 ( .A(_4696__bF_buf1), .B(_3846__bF_buf0), .C(_3856_), .Y(_868_) );
OAI21X1 OAI21X1_3943 ( .A(_4917__bF_buf9), .B(_3844__bF_buf6), .C(cpuregs_19_[10]), .Y(_3857_) );
OAI21X1 OAI21X1_3944 ( .A(_4703__bF_buf1), .B(_3846__bF_buf4), .C(_3857_), .Y(_869_) );
OAI21X1 OAI21X1_3945 ( .A(_4917__bF_buf8), .B(_3844__bF_buf5), .C(cpuregs_19_[11]), .Y(_3858_) );
OAI21X1 OAI21X1_3946 ( .A(_4713__bF_buf1), .B(_3846__bF_buf3), .C(_3858_), .Y(_870_) );
OAI21X1 OAI21X1_3947 ( .A(_4917__bF_buf7), .B(_3844__bF_buf4), .C(cpuregs_19_[12]), .Y(_3859_) );
OAI21X1 OAI21X1_3948 ( .A(_4722__bF_buf1), .B(_3846__bF_buf2), .C(_3859_), .Y(_871_) );
OAI21X1 OAI21X1_3949 ( .A(_4917__bF_buf6), .B(_3844__bF_buf3), .C(cpuregs_19_[13]), .Y(_3860_) );
OAI21X1 OAI21X1_3950 ( .A(_4731__bF_buf1), .B(_3846__bF_buf1), .C(_3860_), .Y(_872_) );
OAI21X1 OAI21X1_3951 ( .A(_4917__bF_buf5), .B(_3844__bF_buf2), .C(cpuregs_19_[14]), .Y(_3861_) );
OAI21X1 OAI21X1_3952 ( .A(_4740__bF_buf1), .B(_3846__bF_buf0), .C(_3861_), .Y(_873_) );
OAI21X1 OAI21X1_3953 ( .A(_4917__bF_buf4), .B(_3844__bF_buf1), .C(cpuregs_19_[15]), .Y(_3862_) );
OAI21X1 OAI21X1_3954 ( .A(_4747__bF_buf1), .B(_3846__bF_buf4), .C(_3862_), .Y(_874_) );
OAI21X1 OAI21X1_3955 ( .A(_4917__bF_buf3), .B(_3844__bF_buf0), .C(cpuregs_19_[16]), .Y(_3863_) );
OAI21X1 OAI21X1_3956 ( .A(_4755__bF_buf1), .B(_3846__bF_buf3), .C(_3863_), .Y(_875_) );
OAI21X1 OAI21X1_3957 ( .A(_4917__bF_buf2), .B(_3844__bF_buf8), .C(cpuregs_19_[17]), .Y(_3864_) );
OAI21X1 OAI21X1_3958 ( .A(_4763__bF_buf1), .B(_3846__bF_buf2), .C(_3864_), .Y(_876_) );
OAI21X1 OAI21X1_3959 ( .A(_4917__bF_buf1), .B(_3844__bF_buf7), .C(cpuregs_19_[18]), .Y(_3865_) );
OAI21X1 OAI21X1_3960 ( .A(_4783__bF_buf1), .B(_3846__bF_buf1), .C(_3865_), .Y(_877_) );
OAI21X1 OAI21X1_3961 ( .A(_4917__bF_buf0), .B(_3844__bF_buf6), .C(cpuregs_19_[19]), .Y(_3866_) );
OAI21X1 OAI21X1_3962 ( .A(_4793__bF_buf1), .B(_3846__bF_buf0), .C(_3866_), .Y(_878_) );
OAI21X1 OAI21X1_3963 ( .A(_4917__bF_buf10), .B(_3844__bF_buf5), .C(cpuregs_19_[20]), .Y(_3867_) );
OAI21X1 OAI21X1_3964 ( .A(_4806__bF_buf1), .B(_3846__bF_buf4), .C(_3867_), .Y(_879_) );
OAI21X1 OAI21X1_3965 ( .A(_4917__bF_buf9), .B(_3844__bF_buf4), .C(cpuregs_19_[21]), .Y(_3868_) );
OAI21X1 OAI21X1_3966 ( .A(_4816__bF_buf1), .B(_3846__bF_buf3), .C(_3868_), .Y(_880_) );
OAI21X1 OAI21X1_3967 ( .A(_4917__bF_buf8), .B(_3844__bF_buf3), .C(cpuregs_19_[22]), .Y(_3869_) );
OAI21X1 OAI21X1_3968 ( .A(_4824__bF_buf1), .B(_3846__bF_buf2), .C(_3869_), .Y(_881_) );
OAI21X1 OAI21X1_3969 ( .A(_4917__bF_buf7), .B(_3844__bF_buf2), .C(cpuregs_19_[23]), .Y(_3870_) );
OAI21X1 OAI21X1_3970 ( .A(_4833__bF_buf1), .B(_3846__bF_buf1), .C(_3870_), .Y(_882_) );
OAI21X1 OAI21X1_3971 ( .A(_4917__bF_buf6), .B(_3844__bF_buf1), .C(cpuregs_19_[24]), .Y(_3871_) );
OAI21X1 OAI21X1_3972 ( .A(_4845__bF_buf1), .B(_3846__bF_buf0), .C(_3871_), .Y(_883_) );
OAI21X1 OAI21X1_3973 ( .A(_4917__bF_buf5), .B(_3844__bF_buf0), .C(cpuregs_19_[25]), .Y(_3872_) );
OAI21X1 OAI21X1_3974 ( .A(_4854__bF_buf1), .B(_3846__bF_buf4), .C(_3872_), .Y(_884_) );
OAI21X1 OAI21X1_3975 ( .A(_4917__bF_buf4), .B(_3844__bF_buf8), .C(cpuregs_19_[26]), .Y(_3873_) );
OAI21X1 OAI21X1_3976 ( .A(_4863__bF_buf1), .B(_3846__bF_buf3), .C(_3873_), .Y(_885_) );
OAI21X1 OAI21X1_3977 ( .A(_4917__bF_buf3), .B(_3844__bF_buf7), .C(cpuregs_19_[27]), .Y(_3874_) );
OAI21X1 OAI21X1_3978 ( .A(_4871__bF_buf1), .B(_3846__bF_buf2), .C(_3874_), .Y(_886_) );
OAI21X1 OAI21X1_3979 ( .A(_4917__bF_buf2), .B(_3844__bF_buf6), .C(cpuregs_19_[28]), .Y(_3875_) );
OAI21X1 OAI21X1_3980 ( .A(_4884__bF_buf1), .B(_3846__bF_buf1), .C(_3875_), .Y(_887_) );
OAI21X1 OAI21X1_3981 ( .A(_4917__bF_buf1), .B(_3844__bF_buf5), .C(cpuregs_19_[29]), .Y(_3876_) );
OAI21X1 OAI21X1_3982 ( .A(_4893__bF_buf1), .B(_3846__bF_buf0), .C(_3876_), .Y(_888_) );
OAI21X1 OAI21X1_3983 ( .A(_4917__bF_buf0), .B(_3844__bF_buf4), .C(cpuregs_19_[30]), .Y(_3877_) );
OAI21X1 OAI21X1_3984 ( .A(_4901__bF_buf1), .B(_3846__bF_buf4), .C(_3877_), .Y(_889_) );
OAI21X1 OAI21X1_3985 ( .A(_4917__bF_buf10), .B(_3844__bF_buf3), .C(cpuregs_19_[31]), .Y(_3878_) );
OAI21X1 OAI21X1_3986 ( .A(_4910__bF_buf1), .B(_3846__bF_buf3), .C(_3878_), .Y(_890_) );
NOR2X1 NOR2X1_1436 ( .A(_4911_), .B(_4635_), .Y(_3879_) );
NAND2X1 NAND2X1_1256 ( .A(_3879_), .B(_5705_), .Y(_3880_) );
NAND2X1 NAND2X1_1257 ( .A(cpuregs_12_[0]), .B(_3880__bF_buf7), .Y(_3881_) );
OAI21X1 OAI21X1_3987 ( .A(_4925__bF_buf1), .B(_3880__bF_buf6), .C(_3881_), .Y(_891_) );
NAND2X1 NAND2X1_1258 ( .A(cpuregs_12_[1]), .B(_3880__bF_buf5), .Y(_3882_) );
OAI21X1 OAI21X1_3988 ( .A(_4933__bF_buf1), .B(_3880__bF_buf4), .C(_3882_), .Y(_892_) );
NAND2X1 NAND2X1_1259 ( .A(cpuregs_12_[2]), .B(_3880__bF_buf3), .Y(_3883_) );
OAI21X1 OAI21X1_3989 ( .A(_4940__bF_buf1), .B(_3880__bF_buf2), .C(_3883_), .Y(_893_) );
NAND2X1 NAND2X1_1260 ( .A(cpuregs_12_[3]), .B(_3880__bF_buf1), .Y(_3884_) );
OAI21X1 OAI21X1_3990 ( .A(_4948__bF_buf1), .B(_3880__bF_buf0), .C(_3884_), .Y(_894_) );
NAND2X1 NAND2X1_1261 ( .A(cpuregs_12_[4]), .B(_3880__bF_buf7), .Y(_3885_) );
OAI21X1 OAI21X1_3991 ( .A(_4955__bF_buf2), .B(_3880__bF_buf6), .C(_3885_), .Y(_895_) );
NAND2X1 NAND2X1_1262 ( .A(cpuregs_12_[5]), .B(_3880__bF_buf5), .Y(_3886_) );
OAI21X1 OAI21X1_3992 ( .A(_4654__bF_buf2), .B(_3880__bF_buf4), .C(_3886_), .Y(_896_) );
NAND2X1 NAND2X1_1263 ( .A(cpuregs_12_[6]), .B(_3880__bF_buf3), .Y(_3887_) );
OAI21X1 OAI21X1_3993 ( .A(_4664__bF_buf2), .B(_3880__bF_buf2), .C(_3887_), .Y(_897_) );
NAND2X1 NAND2X1_1264 ( .A(cpuregs_12_[7]), .B(_3880__bF_buf1), .Y(_3888_) );
OAI21X1 OAI21X1_3994 ( .A(_4677__bF_buf1), .B(_3880__bF_buf0), .C(_3888_), .Y(_898_) );
NAND2X1 NAND2X1_1265 ( .A(cpuregs_12_[8]), .B(_3880__bF_buf7), .Y(_3889_) );
OAI21X1 OAI21X1_3995 ( .A(_4685__bF_buf2), .B(_3880__bF_buf6), .C(_3889_), .Y(_899_) );
NAND2X1 NAND2X1_1266 ( .A(cpuregs_12_[9]), .B(_3880__bF_buf5), .Y(_3890_) );
OAI21X1 OAI21X1_3996 ( .A(_4696__bF_buf0), .B(_3880__bF_buf4), .C(_3890_), .Y(_900_) );
NAND2X1 NAND2X1_1267 ( .A(cpuregs_12_[10]), .B(_3880__bF_buf3), .Y(_3891_) );
OAI21X1 OAI21X1_3997 ( .A(_4703__bF_buf0), .B(_3880__bF_buf2), .C(_3891_), .Y(_901_) );
NAND2X1 NAND2X1_1268 ( .A(cpuregs_12_[11]), .B(_3880__bF_buf1), .Y(_3892_) );
OAI21X1 OAI21X1_3998 ( .A(_4713__bF_buf0), .B(_3880__bF_buf0), .C(_3892_), .Y(_902_) );
NAND2X1 NAND2X1_1269 ( .A(cpuregs_12_[12]), .B(_3880__bF_buf7), .Y(_3893_) );
OAI21X1 OAI21X1_3999 ( .A(_4722__bF_buf0), .B(_3880__bF_buf6), .C(_3893_), .Y(_903_) );
NAND2X1 NAND2X1_1270 ( .A(cpuregs_12_[13]), .B(_3880__bF_buf5), .Y(_3894_) );
OAI21X1 OAI21X1_4000 ( .A(_4731__bF_buf0), .B(_3880__bF_buf4), .C(_3894_), .Y(_904_) );
NAND2X1 NAND2X1_1271 ( .A(cpuregs_12_[14]), .B(_3880__bF_buf3), .Y(_3895_) );
OAI21X1 OAI21X1_4001 ( .A(_4740__bF_buf0), .B(_3880__bF_buf2), .C(_3895_), .Y(_905_) );
NAND2X1 NAND2X1_1272 ( .A(cpuregs_12_[15]), .B(_3880__bF_buf1), .Y(_3896_) );
OAI21X1 OAI21X1_4002 ( .A(_4747__bF_buf0), .B(_3880__bF_buf0), .C(_3896_), .Y(_906_) );
NAND2X1 NAND2X1_1273 ( .A(cpuregs_12_[16]), .B(_3880__bF_buf7), .Y(_3897_) );
OAI21X1 OAI21X1_4003 ( .A(_4755__bF_buf0), .B(_3880__bF_buf6), .C(_3897_), .Y(_907_) );
NAND2X1 NAND2X1_1274 ( .A(cpuregs_12_[17]), .B(_3880__bF_buf5), .Y(_3898_) );
OAI21X1 OAI21X1_4004 ( .A(_4763__bF_buf0), .B(_3880__bF_buf4), .C(_3898_), .Y(_908_) );
NAND2X1 NAND2X1_1275 ( .A(cpuregs_12_[18]), .B(_3880__bF_buf3), .Y(_3899_) );
OAI21X1 OAI21X1_4005 ( .A(_4783__bF_buf0), .B(_3880__bF_buf2), .C(_3899_), .Y(_909_) );
NAND2X1 NAND2X1_1276 ( .A(cpuregs_12_[19]), .B(_3880__bF_buf1), .Y(_3900_) );
OAI21X1 OAI21X1_4006 ( .A(_4793__bF_buf0), .B(_3880__bF_buf0), .C(_3900_), .Y(_910_) );
NAND2X1 NAND2X1_1277 ( .A(cpuregs_12_[20]), .B(_3880__bF_buf7), .Y(_3901_) );
OAI21X1 OAI21X1_4007 ( .A(_4806__bF_buf0), .B(_3880__bF_buf6), .C(_3901_), .Y(_911_) );
NAND2X1 NAND2X1_1278 ( .A(cpuregs_12_[21]), .B(_3880__bF_buf5), .Y(_3902_) );
OAI21X1 OAI21X1_4008 ( .A(_4816__bF_buf0), .B(_3880__bF_buf4), .C(_3902_), .Y(_912_) );
NAND2X1 NAND2X1_1279 ( .A(cpuregs_12_[22]), .B(_3880__bF_buf3), .Y(_3903_) );
OAI21X1 OAI21X1_4009 ( .A(_4824__bF_buf0), .B(_3880__bF_buf2), .C(_3903_), .Y(_913_) );
NAND2X1 NAND2X1_1280 ( .A(cpuregs_12_[23]), .B(_3880__bF_buf1), .Y(_3904_) );
OAI21X1 OAI21X1_4010 ( .A(_4833__bF_buf0), .B(_3880__bF_buf0), .C(_3904_), .Y(_914_) );
NAND2X1 NAND2X1_1281 ( .A(cpuregs_12_[24]), .B(_3880__bF_buf7), .Y(_3905_) );
OAI21X1 OAI21X1_4011 ( .A(_4845__bF_buf0), .B(_3880__bF_buf6), .C(_3905_), .Y(_915_) );
NAND2X1 NAND2X1_1282 ( .A(cpuregs_12_[25]), .B(_3880__bF_buf5), .Y(_3906_) );
OAI21X1 OAI21X1_4012 ( .A(_4854__bF_buf0), .B(_3880__bF_buf4), .C(_3906_), .Y(_916_) );
NAND2X1 NAND2X1_1283 ( .A(cpuregs_12_[26]), .B(_3880__bF_buf3), .Y(_3907_) );
OAI21X1 OAI21X1_4013 ( .A(_4863__bF_buf0), .B(_3880__bF_buf2), .C(_3907_), .Y(_917_) );
NAND2X1 NAND2X1_1284 ( .A(cpuregs_12_[27]), .B(_3880__bF_buf1), .Y(_3908_) );
OAI21X1 OAI21X1_4014 ( .A(_4871__bF_buf0), .B(_3880__bF_buf0), .C(_3908_), .Y(_918_) );
NAND2X1 NAND2X1_1285 ( .A(cpuregs_12_[28]), .B(_3880__bF_buf7), .Y(_3909_) );
OAI21X1 OAI21X1_4015 ( .A(_4884__bF_buf0), .B(_3880__bF_buf6), .C(_3909_), .Y(_919_) );
NAND2X1 NAND2X1_1286 ( .A(cpuregs_12_[29]), .B(_3880__bF_buf5), .Y(_3910_) );
OAI21X1 OAI21X1_4016 ( .A(_4893__bF_buf0), .B(_3880__bF_buf4), .C(_3910_), .Y(_920_) );
NAND2X1 NAND2X1_1287 ( .A(cpuregs_12_[30]), .B(_3880__bF_buf3), .Y(_3911_) );
OAI21X1 OAI21X1_4017 ( .A(_4901__bF_buf0), .B(_3880__bF_buf2), .C(_3911_), .Y(_921_) );
NAND2X1 NAND2X1_1288 ( .A(cpuregs_12_[31]), .B(_3880__bF_buf1), .Y(_3912_) );
OAI21X1 OAI21X1_4018 ( .A(_4910__bF_buf0), .B(_3880__bF_buf0), .C(_3912_), .Y(_922_) );
NOR2X1 NOR2X1_1437 ( .A(_3844__bF_buf2), .B(_5281__bF_buf8), .Y(_3913_) );
INVX1 INVX1_1352 ( .A(_3913_), .Y(_3914_) );
OAI21X1 OAI21X1_4019 ( .A(_5281__bF_buf7), .B(_3844__bF_buf1), .C(cpuregs_18_[0]), .Y(_3915_) );
OAI21X1 OAI21X1_4020 ( .A(_3914__bF_buf4), .B(_4925__bF_buf0), .C(_3915_), .Y(_923_) );
OAI21X1 OAI21X1_4021 ( .A(_5281__bF_buf6), .B(_3844__bF_buf0), .C(cpuregs_18_[1]), .Y(_3916_) );
OAI21X1 OAI21X1_4022 ( .A(_3914__bF_buf3), .B(_4933__bF_buf0), .C(_3916_), .Y(_924_) );
OAI21X1 OAI21X1_4023 ( .A(_5281__bF_buf5), .B(_3844__bF_buf8), .C(cpuregs_18_[2]), .Y(_3917_) );
OAI21X1 OAI21X1_4024 ( .A(_3914__bF_buf2), .B(_4940__bF_buf0), .C(_3917_), .Y(_925_) );
OAI21X1 OAI21X1_4025 ( .A(_5281__bF_buf4), .B(_3844__bF_buf7), .C(cpuregs_18_[3]), .Y(_3918_) );
OAI21X1 OAI21X1_4026 ( .A(_3914__bF_buf1), .B(_4948__bF_buf0), .C(_3918_), .Y(_926_) );
OAI21X1 OAI21X1_4027 ( .A(_5281__bF_buf3), .B(_3844__bF_buf6), .C(cpuregs_18_[4]), .Y(_3919_) );
OAI21X1 OAI21X1_4028 ( .A(_3914__bF_buf0), .B(_4955__bF_buf1), .C(_3919_), .Y(_927_) );
OAI21X1 OAI21X1_4029 ( .A(_5281__bF_buf2), .B(_3844__bF_buf5), .C(cpuregs_18_[5]), .Y(_3920_) );
OAI21X1 OAI21X1_4030 ( .A(_3914__bF_buf4), .B(_4654__bF_buf1), .C(_3920_), .Y(_928_) );
OAI21X1 OAI21X1_4031 ( .A(_5281__bF_buf1), .B(_3844__bF_buf4), .C(cpuregs_18_[6]), .Y(_3921_) );
OAI21X1 OAI21X1_4032 ( .A(_4664__bF_buf1), .B(_3914__bF_buf3), .C(_3921_), .Y(_929_) );
OAI21X1 OAI21X1_4033 ( .A(_5281__bF_buf0), .B(_3844__bF_buf3), .C(cpuregs_18_[7]), .Y(_3922_) );
OAI21X1 OAI21X1_4034 ( .A(_4677__bF_buf0), .B(_3914__bF_buf2), .C(_3922_), .Y(_930_) );
OAI21X1 OAI21X1_4035 ( .A(_5281__bF_buf10), .B(_3844__bF_buf2), .C(cpuregs_18_[8]), .Y(_3923_) );
OAI21X1 OAI21X1_4036 ( .A(_4685__bF_buf1), .B(_3914__bF_buf1), .C(_3923_), .Y(_931_) );
OAI21X1 OAI21X1_4037 ( .A(_5281__bF_buf9), .B(_3844__bF_buf1), .C(cpuregs_18_[9]), .Y(_3924_) );
OAI21X1 OAI21X1_4038 ( .A(_4696__bF_buf4), .B(_3914__bF_buf0), .C(_3924_), .Y(_932_) );
OAI21X1 OAI21X1_4039 ( .A(_5281__bF_buf8), .B(_3844__bF_buf0), .C(cpuregs_18_[10]), .Y(_3925_) );
OAI21X1 OAI21X1_4040 ( .A(_4703__bF_buf4), .B(_3914__bF_buf4), .C(_3925_), .Y(_933_) );
OAI21X1 OAI21X1_4041 ( .A(_5281__bF_buf7), .B(_3844__bF_buf8), .C(cpuregs_18_[11]), .Y(_3926_) );
OAI21X1 OAI21X1_4042 ( .A(_4713__bF_buf4), .B(_3914__bF_buf3), .C(_3926_), .Y(_934_) );
OAI21X1 OAI21X1_4043 ( .A(_5281__bF_buf6), .B(_3844__bF_buf7), .C(cpuregs_18_[12]), .Y(_3927_) );
OAI21X1 OAI21X1_4044 ( .A(_4722__bF_buf4), .B(_3914__bF_buf2), .C(_3927_), .Y(_935_) );
OAI21X1 OAI21X1_4045 ( .A(_5281__bF_buf5), .B(_3844__bF_buf6), .C(cpuregs_18_[13]), .Y(_3928_) );
OAI21X1 OAI21X1_4046 ( .A(_4731__bF_buf4), .B(_3914__bF_buf1), .C(_3928_), .Y(_936_) );
OAI21X1 OAI21X1_4047 ( .A(_5281__bF_buf4), .B(_3844__bF_buf5), .C(cpuregs_18_[14]), .Y(_3929_) );
OAI21X1 OAI21X1_4048 ( .A(_4740__bF_buf4), .B(_3914__bF_buf0), .C(_3929_), .Y(_937_) );
OAI21X1 OAI21X1_4049 ( .A(_5281__bF_buf3), .B(_3844__bF_buf4), .C(cpuregs_18_[15]), .Y(_3930_) );
OAI21X1 OAI21X1_4050 ( .A(_4747__bF_buf4), .B(_3914__bF_buf4), .C(_3930_), .Y(_938_) );
OAI21X1 OAI21X1_4051 ( .A(_5281__bF_buf2), .B(_3844__bF_buf3), .C(cpuregs_18_[16]), .Y(_3931_) );
OAI21X1 OAI21X1_4052 ( .A(_4755__bF_buf4), .B(_3914__bF_buf3), .C(_3931_), .Y(_939_) );
OAI21X1 OAI21X1_4053 ( .A(_5281__bF_buf1), .B(_3844__bF_buf2), .C(cpuregs_18_[17]), .Y(_3932_) );
OAI21X1 OAI21X1_4054 ( .A(_4763__bF_buf4), .B(_3914__bF_buf2), .C(_3932_), .Y(_940_) );
OAI21X1 OAI21X1_4055 ( .A(_5281__bF_buf0), .B(_3844__bF_buf1), .C(cpuregs_18_[18]), .Y(_3933_) );
OAI21X1 OAI21X1_4056 ( .A(_4783__bF_buf4), .B(_3914__bF_buf1), .C(_3933_), .Y(_941_) );
OAI21X1 OAI21X1_4057 ( .A(_5281__bF_buf10), .B(_3844__bF_buf0), .C(cpuregs_18_[19]), .Y(_3934_) );
OAI21X1 OAI21X1_4058 ( .A(_4793__bF_buf4), .B(_3914__bF_buf0), .C(_3934_), .Y(_942_) );
OAI21X1 OAI21X1_4059 ( .A(_5281__bF_buf9), .B(_3844__bF_buf8), .C(cpuregs_18_[20]), .Y(_3935_) );
OAI21X1 OAI21X1_4060 ( .A(_4806__bF_buf4), .B(_3914__bF_buf4), .C(_3935_), .Y(_943_) );
OAI21X1 OAI21X1_4061 ( .A(_5281__bF_buf8), .B(_3844__bF_buf7), .C(cpuregs_18_[21]), .Y(_3936_) );
OAI21X1 OAI21X1_4062 ( .A(_4816__bF_buf4), .B(_3914__bF_buf3), .C(_3936_), .Y(_944_) );
OAI21X1 OAI21X1_4063 ( .A(_5281__bF_buf7), .B(_3844__bF_buf6), .C(cpuregs_18_[22]), .Y(_3937_) );
OAI21X1 OAI21X1_4064 ( .A(_4824__bF_buf4), .B(_3914__bF_buf2), .C(_3937_), .Y(_945_) );
OAI21X1 OAI21X1_4065 ( .A(_5281__bF_buf6), .B(_3844__bF_buf5), .C(cpuregs_18_[23]), .Y(_3938_) );
OAI21X1 OAI21X1_4066 ( .A(_4833__bF_buf4), .B(_3914__bF_buf1), .C(_3938_), .Y(_946_) );
OAI21X1 OAI21X1_4067 ( .A(_5281__bF_buf5), .B(_3844__bF_buf4), .C(cpuregs_18_[24]), .Y(_3939_) );
OAI21X1 OAI21X1_4068 ( .A(_4845__bF_buf4), .B(_3914__bF_buf0), .C(_3939_), .Y(_947_) );
OAI21X1 OAI21X1_4069 ( .A(_5281__bF_buf4), .B(_3844__bF_buf3), .C(cpuregs_18_[25]), .Y(_3940_) );
OAI21X1 OAI21X1_4070 ( .A(_4854__bF_buf4), .B(_3914__bF_buf4), .C(_3940_), .Y(_948_) );
OAI21X1 OAI21X1_4071 ( .A(_5281__bF_buf3), .B(_3844__bF_buf2), .C(cpuregs_18_[26]), .Y(_3941_) );
OAI21X1 OAI21X1_4072 ( .A(_4863__bF_buf4), .B(_3914__bF_buf3), .C(_3941_), .Y(_949_) );
OAI21X1 OAI21X1_4073 ( .A(_5281__bF_buf2), .B(_3844__bF_buf1), .C(cpuregs_18_[27]), .Y(_3942_) );
OAI21X1 OAI21X1_4074 ( .A(_4871__bF_buf4), .B(_3914__bF_buf2), .C(_3942_), .Y(_950_) );
OAI21X1 OAI21X1_4075 ( .A(_5281__bF_buf1), .B(_3844__bF_buf0), .C(cpuregs_18_[28]), .Y(_3943_) );
OAI21X1 OAI21X1_4076 ( .A(_4884__bF_buf4), .B(_3914__bF_buf1), .C(_3943_), .Y(_951_) );
OAI21X1 OAI21X1_4077 ( .A(_5281__bF_buf0), .B(_3844__bF_buf8), .C(cpuregs_18_[29]), .Y(_3944_) );
OAI21X1 OAI21X1_4078 ( .A(_4893__bF_buf4), .B(_3914__bF_buf0), .C(_3944_), .Y(_952_) );
OAI21X1 OAI21X1_4079 ( .A(_5281__bF_buf10), .B(_3844__bF_buf7), .C(cpuregs_18_[30]), .Y(_3945_) );
OAI21X1 OAI21X1_4080 ( .A(_4901__bF_buf4), .B(_3914__bF_buf4), .C(_3945_), .Y(_953_) );
OAI21X1 OAI21X1_4081 ( .A(_5281__bF_buf9), .B(_3844__bF_buf6), .C(cpuregs_18_[31]), .Y(_3946_) );
OAI21X1 OAI21X1_4082 ( .A(_4910__bF_buf4), .B(_3914__bF_buf3), .C(_3946_), .Y(_954_) );
NAND2X1 NAND2X1_1289 ( .A(_3843_), .B(_5313_), .Y(_3947_) );
NAND2X1 NAND2X1_1290 ( .A(cpuregs_17_[0]), .B(_3947__bF_buf7), .Y(_3948_) );
OAI21X1 OAI21X1_4083 ( .A(_4925__bF_buf4), .B(_3947__bF_buf6), .C(_3948_), .Y(_955_) );
NAND2X1 NAND2X1_1291 ( .A(cpuregs_17_[1]), .B(_3947__bF_buf5), .Y(_3949_) );
OAI21X1 OAI21X1_4084 ( .A(_4933__bF_buf4), .B(_3947__bF_buf4), .C(_3949_), .Y(_956_) );
NAND2X1 NAND2X1_1292 ( .A(cpuregs_17_[2]), .B(_3947__bF_buf3), .Y(_3950_) );
OAI21X1 OAI21X1_4085 ( .A(_4940__bF_buf4), .B(_3947__bF_buf2), .C(_3950_), .Y(_957_) );
NAND2X1 NAND2X1_1293 ( .A(cpuregs_17_[3]), .B(_3947__bF_buf1), .Y(_3951_) );
OAI21X1 OAI21X1_4086 ( .A(_4948__bF_buf4), .B(_3947__bF_buf0), .C(_3951_), .Y(_958_) );
NAND2X1 NAND2X1_1294 ( .A(cpuregs_17_[4]), .B(_3947__bF_buf7), .Y(_3952_) );
OAI21X1 OAI21X1_4087 ( .A(_4955__bF_buf0), .B(_3947__bF_buf6), .C(_3952_), .Y(_959_) );
NAND2X1 NAND2X1_1295 ( .A(cpuregs_17_[5]), .B(_3947__bF_buf5), .Y(_3953_) );
OAI21X1 OAI21X1_4088 ( .A(_4654__bF_buf0), .B(_3947__bF_buf4), .C(_3953_), .Y(_960_) );
NAND2X1 NAND2X1_1296 ( .A(cpuregs_17_[6]), .B(_3947__bF_buf3), .Y(_3954_) );
OAI21X1 OAI21X1_4089 ( .A(_4664__bF_buf0), .B(_3947__bF_buf2), .C(_3954_), .Y(_961_) );
NAND2X1 NAND2X1_1297 ( .A(cpuregs_17_[7]), .B(_3947__bF_buf1), .Y(_3955_) );
OAI21X1 OAI21X1_4090 ( .A(_4677__bF_buf4), .B(_3947__bF_buf0), .C(_3955_), .Y(_962_) );
NAND2X1 NAND2X1_1298 ( .A(cpuregs_17_[8]), .B(_3947__bF_buf7), .Y(_3956_) );
OAI21X1 OAI21X1_4091 ( .A(_4685__bF_buf0), .B(_3947__bF_buf6), .C(_3956_), .Y(_963_) );
NAND2X1 NAND2X1_1299 ( .A(cpuregs_17_[9]), .B(_3947__bF_buf5), .Y(_3957_) );
OAI21X1 OAI21X1_4092 ( .A(_4696__bF_buf3), .B(_3947__bF_buf4), .C(_3957_), .Y(_964_) );
NAND2X1 NAND2X1_1300 ( .A(cpuregs_17_[10]), .B(_3947__bF_buf3), .Y(_3958_) );
OAI21X1 OAI21X1_4093 ( .A(_4703__bF_buf3), .B(_3947__bF_buf2), .C(_3958_), .Y(_965_) );
NAND2X1 NAND2X1_1301 ( .A(cpuregs_17_[11]), .B(_3947__bF_buf1), .Y(_3959_) );
OAI21X1 OAI21X1_4094 ( .A(_4713__bF_buf3), .B(_3947__bF_buf0), .C(_3959_), .Y(_966_) );
NAND2X1 NAND2X1_1302 ( .A(cpuregs_17_[12]), .B(_3947__bF_buf7), .Y(_3960_) );
OAI21X1 OAI21X1_4095 ( .A(_4722__bF_buf3), .B(_3947__bF_buf6), .C(_3960_), .Y(_967_) );
NAND2X1 NAND2X1_1303 ( .A(cpuregs_17_[13]), .B(_3947__bF_buf5), .Y(_3961_) );
OAI21X1 OAI21X1_4096 ( .A(_4731__bF_buf3), .B(_3947__bF_buf4), .C(_3961_), .Y(_968_) );
NAND2X1 NAND2X1_1304 ( .A(cpuregs_17_[14]), .B(_3947__bF_buf3), .Y(_3962_) );
OAI21X1 OAI21X1_4097 ( .A(_4740__bF_buf3), .B(_3947__bF_buf2), .C(_3962_), .Y(_969_) );
NAND2X1 NAND2X1_1305 ( .A(cpuregs_17_[15]), .B(_3947__bF_buf1), .Y(_3963_) );
OAI21X1 OAI21X1_4098 ( .A(_4747__bF_buf3), .B(_3947__bF_buf0), .C(_3963_), .Y(_970_) );
NAND2X1 NAND2X1_1306 ( .A(cpuregs_17_[16]), .B(_3947__bF_buf7), .Y(_3964_) );
OAI21X1 OAI21X1_4099 ( .A(_4755__bF_buf3), .B(_3947__bF_buf6), .C(_3964_), .Y(_971_) );
NAND2X1 NAND2X1_1307 ( .A(cpuregs_17_[17]), .B(_3947__bF_buf5), .Y(_3965_) );
OAI21X1 OAI21X1_4100 ( .A(_4763__bF_buf3), .B(_3947__bF_buf4), .C(_3965_), .Y(_972_) );
NAND2X1 NAND2X1_1308 ( .A(cpuregs_17_[18]), .B(_3947__bF_buf3), .Y(_3966_) );
OAI21X1 OAI21X1_4101 ( .A(_4783__bF_buf3), .B(_3947__bF_buf2), .C(_3966_), .Y(_973_) );
NAND2X1 NAND2X1_1309 ( .A(cpuregs_17_[19]), .B(_3947__bF_buf1), .Y(_3967_) );
OAI21X1 OAI21X1_4102 ( .A(_4793__bF_buf3), .B(_3947__bF_buf0), .C(_3967_), .Y(_974_) );
NAND2X1 NAND2X1_1310 ( .A(cpuregs_17_[20]), .B(_3947__bF_buf7), .Y(_3968_) );
OAI21X1 OAI21X1_4103 ( .A(_4806__bF_buf3), .B(_3947__bF_buf6), .C(_3968_), .Y(_975_) );
NAND2X1 NAND2X1_1311 ( .A(cpuregs_17_[21]), .B(_3947__bF_buf5), .Y(_3969_) );
OAI21X1 OAI21X1_4104 ( .A(_4816__bF_buf3), .B(_3947__bF_buf4), .C(_3969_), .Y(_976_) );
NAND2X1 NAND2X1_1312 ( .A(cpuregs_17_[22]), .B(_3947__bF_buf3), .Y(_3970_) );
OAI21X1 OAI21X1_4105 ( .A(_4824__bF_buf3), .B(_3947__bF_buf2), .C(_3970_), .Y(_977_) );
NAND2X1 NAND2X1_1313 ( .A(cpuregs_17_[23]), .B(_3947__bF_buf1), .Y(_3971_) );
OAI21X1 OAI21X1_4106 ( .A(_4833__bF_buf3), .B(_3947__bF_buf0), .C(_3971_), .Y(_978_) );
NAND2X1 NAND2X1_1314 ( .A(cpuregs_17_[24]), .B(_3947__bF_buf7), .Y(_3972_) );
OAI21X1 OAI21X1_4107 ( .A(_4845__bF_buf3), .B(_3947__bF_buf6), .C(_3972_), .Y(_979_) );
NAND2X1 NAND2X1_1315 ( .A(cpuregs_17_[25]), .B(_3947__bF_buf5), .Y(_3973_) );
OAI21X1 OAI21X1_4108 ( .A(_4854__bF_buf3), .B(_3947__bF_buf4), .C(_3973_), .Y(_980_) );
NAND2X1 NAND2X1_1316 ( .A(cpuregs_17_[26]), .B(_3947__bF_buf3), .Y(_3974_) );
OAI21X1 OAI21X1_4109 ( .A(_4863__bF_buf3), .B(_3947__bF_buf2), .C(_3974_), .Y(_981_) );
NAND2X1 NAND2X1_1317 ( .A(cpuregs_17_[27]), .B(_3947__bF_buf1), .Y(_3975_) );
OAI21X1 OAI21X1_4110 ( .A(_4871__bF_buf3), .B(_3947__bF_buf0), .C(_3975_), .Y(_982_) );
NAND2X1 NAND2X1_1318 ( .A(cpuregs_17_[28]), .B(_3947__bF_buf7), .Y(_3976_) );
OAI21X1 OAI21X1_4111 ( .A(_4884__bF_buf3), .B(_3947__bF_buf6), .C(_3976_), .Y(_983_) );
NAND2X1 NAND2X1_1319 ( .A(cpuregs_17_[29]), .B(_3947__bF_buf5), .Y(_3977_) );
OAI21X1 OAI21X1_4112 ( .A(_4893__bF_buf3), .B(_3947__bF_buf4), .C(_3977_), .Y(_984_) );
NAND2X1 NAND2X1_1320 ( .A(cpuregs_17_[30]), .B(_3947__bF_buf3), .Y(_3978_) );
OAI21X1 OAI21X1_4113 ( .A(_4901__bF_buf3), .B(_3947__bF_buf2), .C(_3978_), .Y(_985_) );
NAND2X1 NAND2X1_1321 ( .A(cpuregs_17_[31]), .B(_3947__bF_buf1), .Y(_3979_) );
OAI21X1 OAI21X1_4114 ( .A(_4910__bF_buf3), .B(_3947__bF_buf0), .C(_3979_), .Y(_986_) );
NOR2X1 NOR2X1_1438 ( .A(_3844__bF_buf5), .B(_5706__bF_buf11), .Y(_3980_) );
INVX1 INVX1_1353 ( .A(_3980_), .Y(_3981_) );
OAI21X1 OAI21X1_4115 ( .A(_5706__bF_buf10), .B(_3844__bF_buf4), .C(cpuregs_16_[0]), .Y(_3982_) );
OAI21X1 OAI21X1_4116 ( .A(_3981__bF_buf4), .B(_4925__bF_buf3), .C(_3982_), .Y(_987_) );
OAI21X1 OAI21X1_4117 ( .A(_5706__bF_buf9), .B(_3844__bF_buf3), .C(cpuregs_16_[1]), .Y(_3983_) );
OAI21X1 OAI21X1_4118 ( .A(_3981__bF_buf3), .B(_4933__bF_buf3), .C(_3983_), .Y(_988_) );
OAI21X1 OAI21X1_4119 ( .A(_5706__bF_buf8), .B(_3844__bF_buf2), .C(cpuregs_16_[2]), .Y(_3984_) );
OAI21X1 OAI21X1_4120 ( .A(_3981__bF_buf2), .B(_4940__bF_buf3), .C(_3984_), .Y(_989_) );
OAI21X1 OAI21X1_4121 ( .A(_5706__bF_buf7), .B(_3844__bF_buf1), .C(cpuregs_16_[3]), .Y(_3985_) );
OAI21X1 OAI21X1_4122 ( .A(_3981__bF_buf1), .B(_4948__bF_buf3), .C(_3985_), .Y(_990_) );
OAI21X1 OAI21X1_4123 ( .A(_5706__bF_buf6), .B(_3844__bF_buf0), .C(cpuregs_16_[4]), .Y(_3986_) );
OAI21X1 OAI21X1_4124 ( .A(_3981__bF_buf0), .B(_4955__bF_buf4), .C(_3986_), .Y(_991_) );
OAI21X1 OAI21X1_4125 ( .A(_5706__bF_buf5), .B(_3844__bF_buf8), .C(cpuregs_16_[5]), .Y(_3987_) );
OAI21X1 OAI21X1_4126 ( .A(_3981__bF_buf4), .B(_4654__bF_buf4), .C(_3987_), .Y(_992_) );
OAI21X1 OAI21X1_4127 ( .A(_5706__bF_buf4), .B(_3844__bF_buf7), .C(cpuregs_16_[6]), .Y(_3988_) );
OAI21X1 OAI21X1_4128 ( .A(_3981__bF_buf3), .B(_4664__bF_buf4), .C(_3988_), .Y(_993_) );
OAI21X1 OAI21X1_4129 ( .A(_5706__bF_buf3), .B(_3844__bF_buf6), .C(cpuregs_16_[7]), .Y(_3989_) );
OAI21X1 OAI21X1_4130 ( .A(_3981__bF_buf2), .B(_4677__bF_buf3), .C(_3989_), .Y(_994_) );
OAI21X1 OAI21X1_4131 ( .A(_5706__bF_buf2), .B(_3844__bF_buf5), .C(cpuregs_16_[8]), .Y(_3990_) );
OAI21X1 OAI21X1_4132 ( .A(_4685__bF_buf4), .B(_3981__bF_buf1), .C(_3990_), .Y(_995_) );
OAI21X1 OAI21X1_4133 ( .A(_5706__bF_buf1), .B(_3844__bF_buf4), .C(cpuregs_16_[9]), .Y(_3991_) );
OAI21X1 OAI21X1_4134 ( .A(_4696__bF_buf2), .B(_3981__bF_buf0), .C(_3991_), .Y(_996_) );
OAI21X1 OAI21X1_4135 ( .A(_5706__bF_buf0), .B(_3844__bF_buf3), .C(cpuregs_16_[10]), .Y(_3992_) );
OAI21X1 OAI21X1_4136 ( .A(_4703__bF_buf2), .B(_3981__bF_buf4), .C(_3992_), .Y(_997_) );
OAI21X1 OAI21X1_4137 ( .A(_5706__bF_buf11), .B(_3844__bF_buf2), .C(cpuregs_16_[11]), .Y(_3993_) );
OAI21X1 OAI21X1_4138 ( .A(_4713__bF_buf2), .B(_3981__bF_buf3), .C(_3993_), .Y(_998_) );
OAI21X1 OAI21X1_4139 ( .A(_5706__bF_buf10), .B(_3844__bF_buf1), .C(cpuregs_16_[12]), .Y(_3994_) );
OAI21X1 OAI21X1_4140 ( .A(_4722__bF_buf2), .B(_3981__bF_buf2), .C(_3994_), .Y(_999_) );
OAI21X1 OAI21X1_4141 ( .A(_5706__bF_buf9), .B(_3844__bF_buf0), .C(cpuregs_16_[13]), .Y(_3995_) );
OAI21X1 OAI21X1_4142 ( .A(_4731__bF_buf2), .B(_3981__bF_buf1), .C(_3995_), .Y(_1000_) );
OAI21X1 OAI21X1_4143 ( .A(_5706__bF_buf8), .B(_3844__bF_buf8), .C(cpuregs_16_[14]), .Y(_3996_) );
OAI21X1 OAI21X1_4144 ( .A(_4740__bF_buf2), .B(_3981__bF_buf0), .C(_3996_), .Y(_1001_) );
OAI21X1 OAI21X1_4145 ( .A(_5706__bF_buf7), .B(_3844__bF_buf7), .C(cpuregs_16_[15]), .Y(_3997_) );
OAI21X1 OAI21X1_4146 ( .A(_4747__bF_buf2), .B(_3981__bF_buf4), .C(_3997_), .Y(_1002_) );
OAI21X1 OAI21X1_4147 ( .A(_5706__bF_buf6), .B(_3844__bF_buf6), .C(cpuregs_16_[16]), .Y(_3998_) );
OAI21X1 OAI21X1_4148 ( .A(_4755__bF_buf2), .B(_3981__bF_buf3), .C(_3998_), .Y(_1003_) );
OAI21X1 OAI21X1_4149 ( .A(_5706__bF_buf5), .B(_3844__bF_buf5), .C(cpuregs_16_[17]), .Y(_3999_) );
OAI21X1 OAI21X1_4150 ( .A(_4763__bF_buf2), .B(_3981__bF_buf2), .C(_3999_), .Y(_1004_) );
OAI21X1 OAI21X1_4151 ( .A(_5706__bF_buf4), .B(_3844__bF_buf4), .C(cpuregs_16_[18]), .Y(_4000_) );
OAI21X1 OAI21X1_4152 ( .A(_4783__bF_buf2), .B(_3981__bF_buf1), .C(_4000_), .Y(_1005_) );
OAI21X1 OAI21X1_4153 ( .A(_5706__bF_buf3), .B(_3844__bF_buf3), .C(cpuregs_16_[19]), .Y(_4001_) );
OAI21X1 OAI21X1_4154 ( .A(_4793__bF_buf2), .B(_3981__bF_buf0), .C(_4001_), .Y(_1006_) );
OAI21X1 OAI21X1_4155 ( .A(_5706__bF_buf2), .B(_3844__bF_buf2), .C(cpuregs_16_[20]), .Y(_4002_) );
OAI21X1 OAI21X1_4156 ( .A(_4806__bF_buf2), .B(_3981__bF_buf4), .C(_4002_), .Y(_1007_) );
OAI21X1 OAI21X1_4157 ( .A(_5706__bF_buf1), .B(_3844__bF_buf1), .C(cpuregs_16_[21]), .Y(_4003_) );
OAI21X1 OAI21X1_4158 ( .A(_4816__bF_buf2), .B(_3981__bF_buf3), .C(_4003_), .Y(_1008_) );
OAI21X1 OAI21X1_4159 ( .A(_5706__bF_buf0), .B(_3844__bF_buf0), .C(cpuregs_16_[22]), .Y(_4004_) );
OAI21X1 OAI21X1_4160 ( .A(_4824__bF_buf2), .B(_3981__bF_buf2), .C(_4004_), .Y(_1009_) );
OAI21X1 OAI21X1_4161 ( .A(_5706__bF_buf11), .B(_3844__bF_buf8), .C(cpuregs_16_[23]), .Y(_4005_) );
OAI21X1 OAI21X1_4162 ( .A(_4833__bF_buf2), .B(_3981__bF_buf1), .C(_4005_), .Y(_1010_) );
OAI21X1 OAI21X1_4163 ( .A(_5706__bF_buf10), .B(_3844__bF_buf7), .C(cpuregs_16_[24]), .Y(_4006_) );
OAI21X1 OAI21X1_4164 ( .A(_4845__bF_buf2), .B(_3981__bF_buf0), .C(_4006_), .Y(_1011_) );
OAI21X1 OAI21X1_4165 ( .A(_5706__bF_buf9), .B(_3844__bF_buf6), .C(cpuregs_16_[25]), .Y(_4007_) );
OAI21X1 OAI21X1_4166 ( .A(_4854__bF_buf2), .B(_3981__bF_buf4), .C(_4007_), .Y(_1012_) );
OAI21X1 OAI21X1_4167 ( .A(_5706__bF_buf8), .B(_3844__bF_buf5), .C(cpuregs_16_[26]), .Y(_4008_) );
OAI21X1 OAI21X1_4168 ( .A(_4863__bF_buf2), .B(_3981__bF_buf3), .C(_4008_), .Y(_1013_) );
OAI21X1 OAI21X1_4169 ( .A(_5706__bF_buf7), .B(_3844__bF_buf4), .C(cpuregs_16_[27]), .Y(_4009_) );
OAI21X1 OAI21X1_4170 ( .A(_4871__bF_buf2), .B(_3981__bF_buf2), .C(_4009_), .Y(_1014_) );
OAI21X1 OAI21X1_4171 ( .A(_5706__bF_buf6), .B(_3844__bF_buf3), .C(cpuregs_16_[28]), .Y(_4010_) );
OAI21X1 OAI21X1_4172 ( .A(_4884__bF_buf2), .B(_3981__bF_buf1), .C(_4010_), .Y(_1015_) );
OAI21X1 OAI21X1_4173 ( .A(_5706__bF_buf5), .B(_3844__bF_buf2), .C(cpuregs_16_[29]), .Y(_4011_) );
OAI21X1 OAI21X1_4174 ( .A(_4893__bF_buf2), .B(_3981__bF_buf0), .C(_4011_), .Y(_1016_) );
OAI21X1 OAI21X1_4175 ( .A(_5706__bF_buf4), .B(_3844__bF_buf1), .C(cpuregs_16_[30]), .Y(_4012_) );
OAI21X1 OAI21X1_4176 ( .A(_4901__bF_buf2), .B(_3981__bF_buf4), .C(_4012_), .Y(_1017_) );
OAI21X1 OAI21X1_4177 ( .A(_5706__bF_buf3), .B(_3844__bF_buf0), .C(cpuregs_16_[31]), .Y(_4013_) );
OAI21X1 OAI21X1_4178 ( .A(_4910__bF_buf2), .B(_3981__bF_buf3), .C(_4013_), .Y(_1018_) );
NAND2X1 NAND2X1_1322 ( .A(_3879_), .B(_5745_), .Y(_4014_) );
NAND2X1 NAND2X1_1323 ( .A(cpuregs_15_[0]), .B(_4014__bF_buf7), .Y(_4015_) );
OAI21X1 OAI21X1_4179 ( .A(_4925__bF_buf2), .B(_4014__bF_buf6), .C(_4015_), .Y(_1019_) );
NAND2X1 NAND2X1_1324 ( .A(cpuregs_15_[1]), .B(_4014__bF_buf5), .Y(_4016_) );
OAI21X1 OAI21X1_4180 ( .A(_4933__bF_buf2), .B(_4014__bF_buf4), .C(_4016_), .Y(_1020_) );
NAND2X1 NAND2X1_1325 ( .A(cpuregs_15_[2]), .B(_4014__bF_buf3), .Y(_4017_) );
OAI21X1 OAI21X1_4181 ( .A(_4940__bF_buf2), .B(_4014__bF_buf2), .C(_4017_), .Y(_1021_) );
NAND2X1 NAND2X1_1326 ( .A(cpuregs_15_[3]), .B(_4014__bF_buf1), .Y(_4018_) );
OAI21X1 OAI21X1_4182 ( .A(_4948__bF_buf2), .B(_4014__bF_buf0), .C(_4018_), .Y(_1022_) );
NAND2X1 NAND2X1_1327 ( .A(cpuregs_15_[4]), .B(_4014__bF_buf7), .Y(_4019_) );
OAI21X1 OAI21X1_4183 ( .A(_4955__bF_buf3), .B(_4014__bF_buf6), .C(_4019_), .Y(_1023_) );
NAND2X1 NAND2X1_1328 ( .A(cpuregs_15_[5]), .B(_4014__bF_buf5), .Y(_4020_) );
OAI21X1 OAI21X1_4184 ( .A(_4654__bF_buf3), .B(_4014__bF_buf4), .C(_4020_), .Y(_1024_) );
NAND2X1 NAND2X1_1329 ( .A(cpuregs_15_[6]), .B(_4014__bF_buf3), .Y(_4021_) );
OAI21X1 OAI21X1_4185 ( .A(_4664__bF_buf3), .B(_4014__bF_buf2), .C(_4021_), .Y(_1025_) );
NAND2X1 NAND2X1_1330 ( .A(cpuregs_15_[7]), .B(_4014__bF_buf1), .Y(_4022_) );
OAI21X1 OAI21X1_4186 ( .A(_4677__bF_buf2), .B(_4014__bF_buf0), .C(_4022_), .Y(_1026_) );
NAND2X1 NAND2X1_1331 ( .A(cpuregs_15_[8]), .B(_4014__bF_buf7), .Y(_4023_) );
OAI21X1 OAI21X1_4187 ( .A(_4685__bF_buf3), .B(_4014__bF_buf6), .C(_4023_), .Y(_1027_) );
NAND2X1 NAND2X1_1332 ( .A(cpuregs_15_[9]), .B(_4014__bF_buf5), .Y(_4024_) );
OAI21X1 OAI21X1_4188 ( .A(_4696__bF_buf1), .B(_4014__bF_buf4), .C(_4024_), .Y(_1028_) );
NAND2X1 NAND2X1_1333 ( .A(cpuregs_15_[10]), .B(_4014__bF_buf3), .Y(_4025_) );
OAI21X1 OAI21X1_4189 ( .A(_4703__bF_buf1), .B(_4014__bF_buf2), .C(_4025_), .Y(_1029_) );
NAND2X1 NAND2X1_1334 ( .A(cpuregs_15_[11]), .B(_4014__bF_buf1), .Y(_4026_) );
OAI21X1 OAI21X1_4190 ( .A(_4713__bF_buf1), .B(_4014__bF_buf0), .C(_4026_), .Y(_1030_) );
NAND2X1 NAND2X1_1335 ( .A(cpuregs_15_[12]), .B(_4014__bF_buf7), .Y(_4027_) );
OAI21X1 OAI21X1_4191 ( .A(_4722__bF_buf1), .B(_4014__bF_buf6), .C(_4027_), .Y(_1031_) );
NAND2X1 NAND2X1_1336 ( .A(cpuregs_15_[13]), .B(_4014__bF_buf5), .Y(_4028_) );
OAI21X1 OAI21X1_4192 ( .A(_4731__bF_buf1), .B(_4014__bF_buf4), .C(_4028_), .Y(_1032_) );
NAND2X1 NAND2X1_1337 ( .A(cpuregs_15_[14]), .B(_4014__bF_buf3), .Y(_4029_) );
OAI21X1 OAI21X1_4193 ( .A(_4740__bF_buf1), .B(_4014__bF_buf2), .C(_4029_), .Y(_1033_) );
NAND2X1 NAND2X1_1338 ( .A(cpuregs_15_[15]), .B(_4014__bF_buf1), .Y(_4030_) );
OAI21X1 OAI21X1_4194 ( .A(_4747__bF_buf1), .B(_4014__bF_buf0), .C(_4030_), .Y(_1034_) );
NAND2X1 NAND2X1_1339 ( .A(cpuregs_15_[16]), .B(_4014__bF_buf7), .Y(_4031_) );
OAI21X1 OAI21X1_4195 ( .A(_4755__bF_buf1), .B(_4014__bF_buf6), .C(_4031_), .Y(_1035_) );
NAND2X1 NAND2X1_1340 ( .A(cpuregs_15_[17]), .B(_4014__bF_buf5), .Y(_4032_) );
OAI21X1 OAI21X1_4196 ( .A(_4763__bF_buf1), .B(_4014__bF_buf4), .C(_4032_), .Y(_1036_) );
NAND2X1 NAND2X1_1341 ( .A(cpuregs_15_[18]), .B(_4014__bF_buf3), .Y(_4033_) );
OAI21X1 OAI21X1_4197 ( .A(_4783__bF_buf1), .B(_4014__bF_buf2), .C(_4033_), .Y(_1037_) );
NAND2X1 NAND2X1_1342 ( .A(cpuregs_15_[19]), .B(_4014__bF_buf1), .Y(_4034_) );
OAI21X1 OAI21X1_4198 ( .A(_4793__bF_buf1), .B(_4014__bF_buf0), .C(_4034_), .Y(_1038_) );
NAND2X1 NAND2X1_1343 ( .A(cpuregs_15_[20]), .B(_4014__bF_buf7), .Y(_4035_) );
OAI21X1 OAI21X1_4199 ( .A(_4806__bF_buf1), .B(_4014__bF_buf6), .C(_4035_), .Y(_1039_) );
NAND2X1 NAND2X1_1344 ( .A(cpuregs_15_[21]), .B(_4014__bF_buf5), .Y(_4036_) );
OAI21X1 OAI21X1_4200 ( .A(_4816__bF_buf1), .B(_4014__bF_buf4), .C(_4036_), .Y(_1040_) );
NAND2X1 NAND2X1_1345 ( .A(cpuregs_15_[22]), .B(_4014__bF_buf3), .Y(_4037_) );
OAI21X1 OAI21X1_4201 ( .A(_4824__bF_buf1), .B(_4014__bF_buf2), .C(_4037_), .Y(_1041_) );
NAND2X1 NAND2X1_1346 ( .A(cpuregs_15_[23]), .B(_4014__bF_buf1), .Y(_4038_) );
OAI21X1 OAI21X1_4202 ( .A(_4833__bF_buf1), .B(_4014__bF_buf0), .C(_4038_), .Y(_1042_) );
NAND2X1 NAND2X1_1347 ( .A(cpuregs_15_[24]), .B(_4014__bF_buf7), .Y(_4039_) );
OAI21X1 OAI21X1_4203 ( .A(_4845__bF_buf1), .B(_4014__bF_buf6), .C(_4039_), .Y(_1043_) );
NAND2X1 NAND2X1_1348 ( .A(cpuregs_15_[25]), .B(_4014__bF_buf5), .Y(_4040_) );
OAI21X1 OAI21X1_4204 ( .A(_4854__bF_buf1), .B(_4014__bF_buf4), .C(_4040_), .Y(_1044_) );
NAND2X1 NAND2X1_1349 ( .A(cpuregs_15_[26]), .B(_4014__bF_buf3), .Y(_4041_) );
OAI21X1 OAI21X1_4205 ( .A(_4863__bF_buf1), .B(_4014__bF_buf2), .C(_4041_), .Y(_1045_) );
NAND2X1 NAND2X1_1350 ( .A(cpuregs_15_[27]), .B(_4014__bF_buf1), .Y(_4042_) );
OAI21X1 OAI21X1_4206 ( .A(_4871__bF_buf1), .B(_4014__bF_buf0), .C(_4042_), .Y(_1046_) );
NAND2X1 NAND2X1_1351 ( .A(cpuregs_15_[28]), .B(_4014__bF_buf7), .Y(_4043_) );
OAI21X1 OAI21X1_4207 ( .A(_4884__bF_buf1), .B(_4014__bF_buf6), .C(_4043_), .Y(_1047_) );
NAND2X1 NAND2X1_1352 ( .A(cpuregs_15_[29]), .B(_4014__bF_buf5), .Y(_4044_) );
OAI21X1 OAI21X1_4208 ( .A(_4893__bF_buf1), .B(_4014__bF_buf4), .C(_4044_), .Y(_1048_) );
NAND2X1 NAND2X1_1353 ( .A(cpuregs_15_[30]), .B(_4014__bF_buf3), .Y(_4045_) );
OAI21X1 OAI21X1_4209 ( .A(_4901__bF_buf1), .B(_4014__bF_buf2), .C(_4045_), .Y(_1049_) );
NAND2X1 NAND2X1_1354 ( .A(cpuregs_15_[31]), .B(_4014__bF_buf1), .Y(_4046_) );
OAI21X1 OAI21X1_4210 ( .A(_4910__bF_buf1), .B(_4014__bF_buf0), .C(_4046_), .Y(_1050_) );
NAND2X1 NAND2X1_1355 ( .A(_3879_), .B(_5779_), .Y(_4047_) );
NAND2X1 NAND2X1_1356 ( .A(cpuregs_14_[0]), .B(_4047__bF_buf7), .Y(_4048_) );
OAI21X1 OAI21X1_4211 ( .A(_4925__bF_buf1), .B(_4047__bF_buf6), .C(_4048_), .Y(_1051_) );
NAND2X1 NAND2X1_1357 ( .A(cpuregs_14_[1]), .B(_4047__bF_buf5), .Y(_4049_) );
OAI21X1 OAI21X1_4212 ( .A(_4933__bF_buf1), .B(_4047__bF_buf4), .C(_4049_), .Y(_1052_) );
NAND2X1 NAND2X1_1358 ( .A(cpuregs_14_[2]), .B(_4047__bF_buf3), .Y(_4050_) );
OAI21X1 OAI21X1_4213 ( .A(_4940__bF_buf1), .B(_4047__bF_buf2), .C(_4050_), .Y(_1053_) );
NAND2X1 NAND2X1_1359 ( .A(cpuregs_14_[3]), .B(_4047__bF_buf1), .Y(_4051_) );
OAI21X1 OAI21X1_4214 ( .A(_4948__bF_buf1), .B(_4047__bF_buf0), .C(_4051_), .Y(_1054_) );
NAND2X1 NAND2X1_1360 ( .A(cpuregs_14_[4]), .B(_4047__bF_buf7), .Y(_4052_) );
OAI21X1 OAI21X1_4215 ( .A(_4955__bF_buf2), .B(_4047__bF_buf6), .C(_4052_), .Y(_1055_) );
NAND2X1 NAND2X1_1361 ( .A(cpuregs_14_[5]), .B(_4047__bF_buf5), .Y(_4053_) );
OAI21X1 OAI21X1_4216 ( .A(_4654__bF_buf2), .B(_4047__bF_buf4), .C(_4053_), .Y(_1056_) );
NAND2X1 NAND2X1_1362 ( .A(cpuregs_14_[6]), .B(_4047__bF_buf3), .Y(_4054_) );
OAI21X1 OAI21X1_4217 ( .A(_4664__bF_buf2), .B(_4047__bF_buf2), .C(_4054_), .Y(_1057_) );
NAND2X1 NAND2X1_1363 ( .A(cpuregs_14_[7]), .B(_4047__bF_buf1), .Y(_4055_) );
OAI21X1 OAI21X1_4218 ( .A(_4677__bF_buf1), .B(_4047__bF_buf0), .C(_4055_), .Y(_1058_) );
NAND2X1 NAND2X1_1364 ( .A(cpuregs_14_[8]), .B(_4047__bF_buf7), .Y(_4056_) );
OAI21X1 OAI21X1_4219 ( .A(_4685__bF_buf2), .B(_4047__bF_buf6), .C(_4056_), .Y(_1059_) );
NAND2X1 NAND2X1_1365 ( .A(cpuregs_14_[9]), .B(_4047__bF_buf5), .Y(_4057_) );
OAI21X1 OAI21X1_4220 ( .A(_4696__bF_buf0), .B(_4047__bF_buf4), .C(_4057_), .Y(_1060_) );
NAND2X1 NAND2X1_1366 ( .A(cpuregs_14_[10]), .B(_4047__bF_buf3), .Y(_4058_) );
OAI21X1 OAI21X1_4221 ( .A(_4703__bF_buf0), .B(_4047__bF_buf2), .C(_4058_), .Y(_1061_) );
NAND2X1 NAND2X1_1367 ( .A(cpuregs_14_[11]), .B(_4047__bF_buf1), .Y(_4059_) );
OAI21X1 OAI21X1_4222 ( .A(_4713__bF_buf0), .B(_4047__bF_buf0), .C(_4059_), .Y(_1062_) );
NAND2X1 NAND2X1_1368 ( .A(cpuregs_14_[12]), .B(_4047__bF_buf7), .Y(_4060_) );
OAI21X1 OAI21X1_4223 ( .A(_4722__bF_buf0), .B(_4047__bF_buf6), .C(_4060_), .Y(_1063_) );
NAND2X1 NAND2X1_1369 ( .A(cpuregs_14_[13]), .B(_4047__bF_buf5), .Y(_4061_) );
OAI21X1 OAI21X1_4224 ( .A(_4731__bF_buf0), .B(_4047__bF_buf4), .C(_4061_), .Y(_1064_) );
NAND2X1 NAND2X1_1370 ( .A(cpuregs_14_[14]), .B(_4047__bF_buf3), .Y(_4062_) );
OAI21X1 OAI21X1_4225 ( .A(_4740__bF_buf0), .B(_4047__bF_buf2), .C(_4062_), .Y(_1065_) );
NAND2X1 NAND2X1_1371 ( .A(cpuregs_14_[15]), .B(_4047__bF_buf1), .Y(_4063_) );
OAI21X1 OAI21X1_4226 ( .A(_4747__bF_buf0), .B(_4047__bF_buf0), .C(_4063_), .Y(_1066_) );
NAND2X1 NAND2X1_1372 ( .A(cpuregs_14_[16]), .B(_4047__bF_buf7), .Y(_4064_) );
OAI21X1 OAI21X1_4227 ( .A(_4755__bF_buf0), .B(_4047__bF_buf6), .C(_4064_), .Y(_1067_) );
NAND2X1 NAND2X1_1373 ( .A(cpuregs_14_[17]), .B(_4047__bF_buf5), .Y(_4065_) );
OAI21X1 OAI21X1_4228 ( .A(_4763__bF_buf0), .B(_4047__bF_buf4), .C(_4065_), .Y(_1068_) );
NAND2X1 NAND2X1_1374 ( .A(cpuregs_14_[18]), .B(_4047__bF_buf3), .Y(_4066_) );
OAI21X1 OAI21X1_4229 ( .A(_4783__bF_buf0), .B(_4047__bF_buf2), .C(_4066_), .Y(_1069_) );
NAND2X1 NAND2X1_1375 ( .A(cpuregs_14_[19]), .B(_4047__bF_buf1), .Y(_4067_) );
OAI21X1 OAI21X1_4230 ( .A(_4793__bF_buf0), .B(_4047__bF_buf0), .C(_4067_), .Y(_1070_) );
NAND2X1 NAND2X1_1376 ( .A(cpuregs_14_[20]), .B(_4047__bF_buf7), .Y(_4068_) );
OAI21X1 OAI21X1_4231 ( .A(_4806__bF_buf0), .B(_4047__bF_buf6), .C(_4068_), .Y(_1071_) );
NAND2X1 NAND2X1_1377 ( .A(cpuregs_14_[21]), .B(_4047__bF_buf5), .Y(_4069_) );
OAI21X1 OAI21X1_4232 ( .A(_4816__bF_buf0), .B(_4047__bF_buf4), .C(_4069_), .Y(_1072_) );
NAND2X1 NAND2X1_1378 ( .A(cpuregs_14_[22]), .B(_4047__bF_buf3), .Y(_4070_) );
OAI21X1 OAI21X1_4233 ( .A(_4824__bF_buf0), .B(_4047__bF_buf2), .C(_4070_), .Y(_1073_) );
NAND2X1 NAND2X1_1379 ( .A(cpuregs_14_[23]), .B(_4047__bF_buf1), .Y(_4071_) );
OAI21X1 OAI21X1_4234 ( .A(_4833__bF_buf0), .B(_4047__bF_buf0), .C(_4071_), .Y(_1074_) );
NAND2X1 NAND2X1_1380 ( .A(cpuregs_14_[24]), .B(_4047__bF_buf7), .Y(_4072_) );
OAI21X1 OAI21X1_4235 ( .A(_4845__bF_buf0), .B(_4047__bF_buf6), .C(_4072_), .Y(_1075_) );
NAND2X1 NAND2X1_1381 ( .A(cpuregs_14_[25]), .B(_4047__bF_buf5), .Y(_4073_) );
OAI21X1 OAI21X1_4236 ( .A(_4854__bF_buf0), .B(_4047__bF_buf4), .C(_4073_), .Y(_1076_) );
NAND2X1 NAND2X1_1382 ( .A(cpuregs_14_[26]), .B(_4047__bF_buf3), .Y(_4074_) );
OAI21X1 OAI21X1_4237 ( .A(_4863__bF_buf0), .B(_4047__bF_buf2), .C(_4074_), .Y(_1077_) );
NAND2X1 NAND2X1_1383 ( .A(cpuregs_14_[27]), .B(_4047__bF_buf1), .Y(_4075_) );
OAI21X1 OAI21X1_4238 ( .A(_4871__bF_buf0), .B(_4047__bF_buf0), .C(_4075_), .Y(_1078_) );
NAND2X1 NAND2X1_1384 ( .A(cpuregs_14_[28]), .B(_4047__bF_buf7), .Y(_4076_) );
OAI21X1 OAI21X1_4239 ( .A(_4884__bF_buf0), .B(_4047__bF_buf6), .C(_4076_), .Y(_1079_) );
NAND2X1 NAND2X1_1385 ( .A(cpuregs_14_[29]), .B(_4047__bF_buf5), .Y(_4077_) );
OAI21X1 OAI21X1_4240 ( .A(_4893__bF_buf0), .B(_4047__bF_buf4), .C(_4077_), .Y(_1080_) );
NAND2X1 NAND2X1_1386 ( .A(cpuregs_14_[30]), .B(_4047__bF_buf3), .Y(_4078_) );
OAI21X1 OAI21X1_4241 ( .A(_4901__bF_buf0), .B(_4047__bF_buf2), .C(_4078_), .Y(_1081_) );
NAND2X1 NAND2X1_1387 ( .A(cpuregs_14_[31]), .B(_4047__bF_buf1), .Y(_4079_) );
OAI21X1 OAI21X1_4242 ( .A(_4910__bF_buf0), .B(_4047__bF_buf0), .C(_4079_), .Y(_1082_) );
NAND2X1 NAND2X1_1388 ( .A(_3879_), .B(_5313_), .Y(_4080_) );
NAND2X1 NAND2X1_1389 ( .A(cpuregs_13_[0]), .B(_4080__bF_buf7), .Y(_4081_) );
OAI21X1 OAI21X1_4243 ( .A(_4925__bF_buf0), .B(_4080__bF_buf6), .C(_4081_), .Y(_1083_) );
NAND2X1 NAND2X1_1390 ( .A(cpuregs_13_[1]), .B(_4080__bF_buf5), .Y(_4082_) );
OAI21X1 OAI21X1_4244 ( .A(_4933__bF_buf0), .B(_4080__bF_buf4), .C(_4082_), .Y(_1084_) );
NAND2X1 NAND2X1_1391 ( .A(cpuregs_13_[2]), .B(_4080__bF_buf3), .Y(_4083_) );
OAI21X1 OAI21X1_4245 ( .A(_4940__bF_buf0), .B(_4080__bF_buf2), .C(_4083_), .Y(_1085_) );
NAND2X1 NAND2X1_1392 ( .A(cpuregs_13_[3]), .B(_4080__bF_buf1), .Y(_4084_) );
OAI21X1 OAI21X1_4246 ( .A(_4948__bF_buf0), .B(_4080__bF_buf0), .C(_4084_), .Y(_1086_) );
NAND2X1 NAND2X1_1393 ( .A(cpuregs_13_[4]), .B(_4080__bF_buf7), .Y(_4085_) );
OAI21X1 OAI21X1_4247 ( .A(_4955__bF_buf1), .B(_4080__bF_buf6), .C(_4085_), .Y(_1087_) );
NAND2X1 NAND2X1_1394 ( .A(cpuregs_13_[5]), .B(_4080__bF_buf5), .Y(_4086_) );
OAI21X1 OAI21X1_4248 ( .A(_4654__bF_buf1), .B(_4080__bF_buf4), .C(_4086_), .Y(_1088_) );
NAND2X1 NAND2X1_1395 ( .A(cpuregs_13_[6]), .B(_4080__bF_buf3), .Y(_4087_) );
OAI21X1 OAI21X1_4249 ( .A(_4664__bF_buf1), .B(_4080__bF_buf2), .C(_4087_), .Y(_1089_) );
NAND2X1 NAND2X1_1396 ( .A(cpuregs_13_[7]), .B(_4080__bF_buf1), .Y(_4088_) );
OAI21X1 OAI21X1_4250 ( .A(_4677__bF_buf0), .B(_4080__bF_buf0), .C(_4088_), .Y(_1090_) );
NAND2X1 NAND2X1_1397 ( .A(cpuregs_13_[8]), .B(_4080__bF_buf7), .Y(_4089_) );
OAI21X1 OAI21X1_4251 ( .A(_4685__bF_buf1), .B(_4080__bF_buf6), .C(_4089_), .Y(_1091_) );
NAND2X1 NAND2X1_1398 ( .A(cpuregs_13_[9]), .B(_4080__bF_buf5), .Y(_4090_) );
OAI21X1 OAI21X1_4252 ( .A(_4696__bF_buf4), .B(_4080__bF_buf4), .C(_4090_), .Y(_1092_) );
NAND2X1 NAND2X1_1399 ( .A(cpuregs_13_[10]), .B(_4080__bF_buf3), .Y(_4091_) );
OAI21X1 OAI21X1_4253 ( .A(_4703__bF_buf4), .B(_4080__bF_buf2), .C(_4091_), .Y(_1093_) );
NAND2X1 NAND2X1_1400 ( .A(cpuregs_13_[11]), .B(_4080__bF_buf1), .Y(_4092_) );
OAI21X1 OAI21X1_4254 ( .A(_4713__bF_buf4), .B(_4080__bF_buf0), .C(_4092_), .Y(_1094_) );
NAND2X1 NAND2X1_1401 ( .A(cpuregs_13_[12]), .B(_4080__bF_buf7), .Y(_4093_) );
OAI21X1 OAI21X1_4255 ( .A(_4722__bF_buf4), .B(_4080__bF_buf6), .C(_4093_), .Y(_1095_) );
NAND2X1 NAND2X1_1402 ( .A(cpuregs_13_[13]), .B(_4080__bF_buf5), .Y(_4094_) );
OAI21X1 OAI21X1_4256 ( .A(_4731__bF_buf4), .B(_4080__bF_buf4), .C(_4094_), .Y(_1096_) );
NAND2X1 NAND2X1_1403 ( .A(cpuregs_13_[14]), .B(_4080__bF_buf3), .Y(_4095_) );
OAI21X1 OAI21X1_4257 ( .A(_4740__bF_buf4), .B(_4080__bF_buf2), .C(_4095_), .Y(_1097_) );
NAND2X1 NAND2X1_1404 ( .A(cpuregs_13_[15]), .B(_4080__bF_buf1), .Y(_4096_) );
OAI21X1 OAI21X1_4258 ( .A(_4747__bF_buf4), .B(_4080__bF_buf0), .C(_4096_), .Y(_1098_) );
NAND2X1 NAND2X1_1405 ( .A(cpuregs_13_[16]), .B(_4080__bF_buf7), .Y(_4097_) );
OAI21X1 OAI21X1_4259 ( .A(_4755__bF_buf4), .B(_4080__bF_buf6), .C(_4097_), .Y(_1099_) );
NAND2X1 NAND2X1_1406 ( .A(cpuregs_13_[17]), .B(_4080__bF_buf5), .Y(_4098_) );
OAI21X1 OAI21X1_4260 ( .A(_4763__bF_buf4), .B(_4080__bF_buf4), .C(_4098_), .Y(_1100_) );
NAND2X1 NAND2X1_1407 ( .A(cpuregs_13_[18]), .B(_4080__bF_buf3), .Y(_4099_) );
OAI21X1 OAI21X1_4261 ( .A(_4783__bF_buf4), .B(_4080__bF_buf2), .C(_4099_), .Y(_1101_) );
NAND2X1 NAND2X1_1408 ( .A(cpuregs_13_[19]), .B(_4080__bF_buf1), .Y(_4100_) );
OAI21X1 OAI21X1_4262 ( .A(_4793__bF_buf4), .B(_4080__bF_buf0), .C(_4100_), .Y(_1102_) );
NAND2X1 NAND2X1_1409 ( .A(cpuregs_13_[20]), .B(_4080__bF_buf7), .Y(_4101_) );
OAI21X1 OAI21X1_4263 ( .A(_4806__bF_buf4), .B(_4080__bF_buf6), .C(_4101_), .Y(_1103_) );
NAND2X1 NAND2X1_1410 ( .A(cpuregs_13_[21]), .B(_4080__bF_buf5), .Y(_4102_) );
OAI21X1 OAI21X1_4264 ( .A(_4816__bF_buf4), .B(_4080__bF_buf4), .C(_4102_), .Y(_1104_) );
NAND2X1 NAND2X1_1411 ( .A(cpuregs_13_[22]), .B(_4080__bF_buf3), .Y(_4103_) );
OAI21X1 OAI21X1_4265 ( .A(_4824__bF_buf4), .B(_4080__bF_buf2), .C(_4103_), .Y(_1105_) );
NAND2X1 NAND2X1_1412 ( .A(cpuregs_13_[23]), .B(_4080__bF_buf1), .Y(_4104_) );
OAI21X1 OAI21X1_4266 ( .A(_4833__bF_buf4), .B(_4080__bF_buf0), .C(_4104_), .Y(_1106_) );
NAND2X1 NAND2X1_1413 ( .A(cpuregs_13_[24]), .B(_4080__bF_buf7), .Y(_4105_) );
OAI21X1 OAI21X1_4267 ( .A(_4845__bF_buf4), .B(_4080__bF_buf6), .C(_4105_), .Y(_1107_) );
NAND2X1 NAND2X1_1414 ( .A(cpuregs_13_[25]), .B(_4080__bF_buf5), .Y(_4106_) );
OAI21X1 OAI21X1_4268 ( .A(_4854__bF_buf4), .B(_4080__bF_buf4), .C(_4106_), .Y(_1108_) );
NAND2X1 NAND2X1_1415 ( .A(cpuregs_13_[26]), .B(_4080__bF_buf3), .Y(_4107_) );
OAI21X1 OAI21X1_4269 ( .A(_4863__bF_buf4), .B(_4080__bF_buf2), .C(_4107_), .Y(_1109_) );
NAND2X1 NAND2X1_1416 ( .A(cpuregs_13_[27]), .B(_4080__bF_buf1), .Y(_4108_) );
OAI21X1 OAI21X1_4270 ( .A(_4871__bF_buf4), .B(_4080__bF_buf0), .C(_4108_), .Y(_1110_) );
NAND2X1 NAND2X1_1417 ( .A(cpuregs_13_[28]), .B(_4080__bF_buf7), .Y(_4109_) );
OAI21X1 OAI21X1_4271 ( .A(_4884__bF_buf4), .B(_4080__bF_buf6), .C(_4109_), .Y(_1111_) );
NAND2X1 NAND2X1_1418 ( .A(cpuregs_13_[29]), .B(_4080__bF_buf5), .Y(_4110_) );
OAI21X1 OAI21X1_4272 ( .A(_4893__bF_buf4), .B(_4080__bF_buf4), .C(_4110_), .Y(_1112_) );
NAND2X1 NAND2X1_1419 ( .A(cpuregs_13_[30]), .B(_4080__bF_buf3), .Y(_4111_) );
OAI21X1 OAI21X1_4273 ( .A(_4901__bF_buf4), .B(_4080__bF_buf2), .C(_4111_), .Y(_1113_) );
NAND2X1 NAND2X1_1420 ( .A(cpuregs_13_[31]), .B(_4080__bF_buf1), .Y(_4112_) );
OAI21X1 OAI21X1_4274 ( .A(_4910__bF_buf4), .B(_4080__bF_buf0), .C(_4112_), .Y(_1114_) );
NOR2X1 NOR2X1_1439 ( .A(count_cycle_0_), .B(_4426__bF_buf10), .Y(_0__0_) );
AND2X2 AND2X2_270 ( .A(count_cycle_0_), .B(count_cycle_1_), .Y(_4113_) );
OAI21X1 OAI21X1_4275 ( .A(count_cycle_0_), .B(count_cycle_1_), .C(resetn_bF_buf0), .Y(_4114_) );
NOR2X1 NOR2X1_1440 ( .A(_4114_), .B(_4113_), .Y(_0__1_) );
NAND2X1 NAND2X1_1421 ( .A(count_cycle_2_), .B(_4113_), .Y(_4115_) );
INVX1 INVX1_1354 ( .A(_4115_), .Y(_4116_) );
OAI21X1 OAI21X1_4276 ( .A(_4113_), .B(count_cycle_2_), .C(resetn_bF_buf11), .Y(_4117_) );
NOR2X1 NOR2X1_1441 ( .A(_4117_), .B(_4116_), .Y(_0__2_) );
INVX1 INVX1_1355 ( .A(count_cycle_3_), .Y(_4118_) );
NOR2X1 NOR2X1_1442 ( .A(_4118_), .B(_4115_), .Y(_4119_) );
OAI21X1 OAI21X1_4277 ( .A(_4116_), .B(count_cycle_3_), .C(resetn_bF_buf10), .Y(_4120_) );
NOR2X1 NOR2X1_1443 ( .A(_4119_), .B(_4120_), .Y(_0__3_) );
AND2X2 AND2X2_271 ( .A(_4119_), .B(count_cycle_4_), .Y(_4121_) );
OAI21X1 OAI21X1_4278 ( .A(_4119_), .B(count_cycle_4_), .C(resetn_bF_buf9), .Y(_4122_) );
NOR2X1 NOR2X1_1444 ( .A(_4122_), .B(_4121_), .Y(_0__4_) );
AND2X2 AND2X2_272 ( .A(_4121_), .B(count_cycle_5_), .Y(_4123_) );
OAI21X1 OAI21X1_4279 ( .A(_4121_), .B(count_cycle_5_), .C(resetn_bF_buf8), .Y(_4124_) );
NOR2X1 NOR2X1_1445 ( .A(_4124_), .B(_4123_), .Y(_0__5_) );
NAND2X1 NAND2X1_1422 ( .A(count_cycle_6_), .B(_4123_), .Y(_4125_) );
INVX1 INVX1_1356 ( .A(_4125_), .Y(_4126_) );
OAI21X1 OAI21X1_4280 ( .A(_4123_), .B(count_cycle_6_), .C(resetn_bF_buf7), .Y(_4127_) );
NOR2X1 NOR2X1_1446 ( .A(_4127_), .B(_4126_), .Y(_0__6_) );
INVX1 INVX1_1357 ( .A(count_cycle_7_), .Y(_4128_) );
NOR2X1 NOR2X1_1447 ( .A(_4128_), .B(_4125_), .Y(_4129_) );
OAI21X1 OAI21X1_4281 ( .A(_4126_), .B(count_cycle_7_), .C(resetn_bF_buf6), .Y(_4130_) );
NOR2X1 NOR2X1_1448 ( .A(_4129_), .B(_4130_), .Y(_0__7_) );
AND2X2 AND2X2_273 ( .A(_4129_), .B(count_cycle_8_), .Y(_4131_) );
OAI21X1 OAI21X1_4282 ( .A(_4129_), .B(count_cycle_8_), .C(resetn_bF_buf5), .Y(_4132_) );
NOR2X1 NOR2X1_1449 ( .A(_4132_), .B(_4131_), .Y(_0__8_) );
AND2X2 AND2X2_274 ( .A(_4131_), .B(count_cycle_9_), .Y(_4133_) );
OAI21X1 OAI21X1_4283 ( .A(_4131_), .B(count_cycle_9_), .C(resetn_bF_buf4), .Y(_4134_) );
NOR2X1 NOR2X1_1450 ( .A(_4134_), .B(_4133_), .Y(_0__9_) );
NAND2X1 NAND2X1_1423 ( .A(count_cycle_10_), .B(_4133_), .Y(_4135_) );
INVX1 INVX1_1358 ( .A(_4135_), .Y(_4136_) );
OAI21X1 OAI21X1_4284 ( .A(_4133_), .B(count_cycle_10_), .C(resetn_bF_buf3), .Y(_4137_) );
NOR2X1 NOR2X1_1451 ( .A(_4137_), .B(_4136_), .Y(_0__10_) );
INVX1 INVX1_1359 ( .A(count_cycle_11_), .Y(_4138_) );
NOR2X1 NOR2X1_1452 ( .A(_4138_), .B(_4135_), .Y(_4139_) );
OAI21X1 OAI21X1_4285 ( .A(_4136_), .B(count_cycle_11_), .C(resetn_bF_buf2), .Y(_4140_) );
NOR2X1 NOR2X1_1453 ( .A(_4139_), .B(_4140_), .Y(_0__11_) );
NAND2X1 NAND2X1_1424 ( .A(count_cycle_12_), .B(_4139_), .Y(_4141_) );
INVX1 INVX1_1360 ( .A(_4141_), .Y(_4142_) );
OAI21X1 OAI21X1_4286 ( .A(_4139_), .B(count_cycle_12_), .C(resetn_bF_buf1), .Y(_4143_) );
NOR2X1 NOR2X1_1454 ( .A(_4143_), .B(_4142_), .Y(_0__12_) );
INVX1 INVX1_1361 ( .A(count_cycle_13_), .Y(_4144_) );
NOR2X1 NOR2X1_1455 ( .A(_4144_), .B(_4141_), .Y(_4145_) );
OAI21X1 OAI21X1_4287 ( .A(_4142_), .B(count_cycle_13_), .C(resetn_bF_buf0), .Y(_4146_) );
NOR2X1 NOR2X1_1456 ( .A(_4145_), .B(_4146_), .Y(_0__13_) );
NAND2X1 NAND2X1_1425 ( .A(count_cycle_14_), .B(_4145_), .Y(_4147_) );
INVX1 INVX1_1362 ( .A(_4147_), .Y(_4148_) );
OAI21X1 OAI21X1_4288 ( .A(_4145_), .B(count_cycle_14_), .C(resetn_bF_buf11), .Y(_4149_) );
NOR2X1 NOR2X1_1457 ( .A(_4149_), .B(_4148_), .Y(_0__14_) );
INVX1 INVX1_1363 ( .A(count_cycle_15_), .Y(_4150_) );
NOR2X1 NOR2X1_1458 ( .A(_4150_), .B(_4147_), .Y(_4151_) );
OAI21X1 OAI21X1_4289 ( .A(_4148_), .B(count_cycle_15_), .C(resetn_bF_buf10), .Y(_4152_) );
NOR2X1 NOR2X1_1459 ( .A(_4151_), .B(_4152_), .Y(_0__15_) );
OAI21X1 OAI21X1_4290 ( .A(_4151_), .B(count_cycle_16_), .C(resetn_bF_buf9), .Y(_4153_) );
AOI21X1 AOI21X1_1062 ( .A(count_cycle_16_), .B(_4151_), .C(_4153_), .Y(_0__16_) );
AOI21X1 AOI21X1_1063 ( .A(count_cycle_16_), .B(_4151_), .C(count_cycle_17_), .Y(_4154_) );
NAND2X1 NAND2X1_1426 ( .A(count_cycle_8_), .B(count_cycle_9_), .Y(_4155_) );
NAND2X1 NAND2X1_1427 ( .A(count_cycle_10_), .B(count_cycle_11_), .Y(_4156_) );
NOR2X1 NOR2X1_1460 ( .A(_4155_), .B(_4156_), .Y(_4157_) );
NAND2X1 NAND2X1_1428 ( .A(count_cycle_12_), .B(count_cycle_13_), .Y(_4158_) );
NAND2X1 NAND2X1_1429 ( .A(count_cycle_14_), .B(count_cycle_15_), .Y(_4159_) );
NOR2X1 NOR2X1_1461 ( .A(_4158_), .B(_4159_), .Y(_4160_) );
NAND2X1 NAND2X1_1430 ( .A(_4157_), .B(_4160_), .Y(_4161_) );
INVX1 INVX1_1364 ( .A(_4161_), .Y(_4162_) );
NAND2X1 NAND2X1_1431 ( .A(_4162_), .B(_4129_), .Y(_4163_) );
NAND2X1 NAND2X1_1432 ( .A(count_cycle_16_), .B(count_cycle_17_), .Y(_4164_) );
OAI21X1 OAI21X1_4291 ( .A(_4163_), .B(_4164_), .C(resetn_bF_buf8), .Y(_4165_) );
NOR2X1 NOR2X1_1462 ( .A(_4165_), .B(_4154_), .Y(_0__17_) );
NOR2X1 NOR2X1_1463 ( .A(_4164_), .B(_4163_), .Y(_4166_) );
AND2X2 AND2X2_275 ( .A(_4166_), .B(count_cycle_18_), .Y(_4167_) );
OAI21X1 OAI21X1_4292 ( .A(_4166_), .B(count_cycle_18_), .C(resetn_bF_buf7), .Y(_4168_) );
NOR2X1 NOR2X1_1464 ( .A(_4168_), .B(_4167_), .Y(_0__18_) );
INVX1 INVX1_1365 ( .A(_4164_), .Y(_4169_) );
NAND3X1 NAND3X1_115 ( .A(count_cycle_18_), .B(count_cycle_19_), .C(_4169_), .Y(_4170_) );
NOR2X1 NOR2X1_1465 ( .A(_4170_), .B(_4163_), .Y(_4171_) );
OAI21X1 OAI21X1_4293 ( .A(_4167_), .B(count_cycle_19_), .C(resetn_bF_buf6), .Y(_4172_) );
NOR2X1 NOR2X1_1466 ( .A(_4171_), .B(_4172_), .Y(_0__19_) );
INVX1 INVX1_1366 ( .A(count_cycle_20_), .Y(_4173_) );
INVX1 INVX1_1367 ( .A(_4171_), .Y(_4174_) );
NOR2X1 NOR2X1_1467 ( .A(_4173_), .B(_4174_), .Y(_4175_) );
OAI21X1 OAI21X1_4294 ( .A(_4171_), .B(count_cycle_20_), .C(resetn_bF_buf5), .Y(_4176_) );
NOR2X1 NOR2X1_1468 ( .A(_4176_), .B(_4175_), .Y(_0__20_) );
INVX1 INVX1_1368 ( .A(count_cycle_21_), .Y(_4177_) );
INVX1 INVX1_1369 ( .A(_4175_), .Y(_4178_) );
NOR2X1 NOR2X1_1469 ( .A(_4173_), .B(_4177_), .Y(_4179_) );
INVX1 INVX1_1370 ( .A(_4179_), .Y(_4180_) );
OAI21X1 OAI21X1_4295 ( .A(_4174_), .B(_4180_), .C(resetn_bF_buf4), .Y(_4181_) );
AOI21X1 AOI21X1_1064 ( .A(_4177_), .B(_4178_), .C(_4181_), .Y(_0__21_) );
NAND2X1 NAND2X1_1433 ( .A(_4179_), .B(_4171_), .Y(_4182_) );
INVX1 INVX1_1371 ( .A(_4182_), .Y(_4183_) );
OAI21X1 OAI21X1_4296 ( .A(_4183_), .B(count_cycle_22_), .C(resetn_bF_buf3), .Y(_4184_) );
AOI21X1 AOI21X1_1065 ( .A(count_cycle_22_), .B(_4183_), .C(_4184_), .Y(_0__22_) );
AOI21X1 AOI21X1_1066 ( .A(count_cycle_22_), .B(_4183_), .C(count_cycle_23_), .Y(_4185_) );
NAND2X1 NAND2X1_1434 ( .A(count_cycle_22_), .B(count_cycle_23_), .Y(_4186_) );
OAI21X1 OAI21X1_4297 ( .A(_4182_), .B(_4186_), .C(resetn_bF_buf2), .Y(_4187_) );
NOR2X1 NOR2X1_1470 ( .A(_4187_), .B(_4185_), .Y(_0__23_) );
INVX1 INVX1_1372 ( .A(count_cycle_24_), .Y(_4188_) );
NOR2X1 NOR2X1_1471 ( .A(_4186_), .B(_4182_), .Y(_4189_) );
INVX1 INVX1_1373 ( .A(_4189_), .Y(_4190_) );
NOR2X1 NOR2X1_1472 ( .A(_4188_), .B(_4190_), .Y(_4191_) );
OAI21X1 OAI21X1_4298 ( .A(_4189_), .B(count_cycle_24_), .C(resetn_bF_buf1), .Y(_4192_) );
NOR2X1 NOR2X1_1473 ( .A(_4192_), .B(_4191_), .Y(_0__24_) );
INVX1 INVX1_1374 ( .A(count_cycle_25_), .Y(_4193_) );
INVX1 INVX1_1375 ( .A(_4191_), .Y(_4194_) );
NOR2X1 NOR2X1_1474 ( .A(_4188_), .B(_4193_), .Y(_4195_) );
INVX1 INVX1_1376 ( .A(_4195_), .Y(_4196_) );
OAI21X1 OAI21X1_4299 ( .A(_4190_), .B(_4196_), .C(resetn_bF_buf0), .Y(_4197_) );
AOI21X1 AOI21X1_1067 ( .A(_4193_), .B(_4194_), .C(_4197_), .Y(_0__25_) );
NAND2X1 NAND2X1_1435 ( .A(_4195_), .B(_4189_), .Y(_4198_) );
INVX1 INVX1_1377 ( .A(_4198_), .Y(_4199_) );
OAI21X1 OAI21X1_4300 ( .A(_4199_), .B(count_cycle_26_), .C(resetn_bF_buf11), .Y(_4200_) );
INVX1 INVX1_1378 ( .A(count_cycle_26_), .Y(_4201_) );
NOR2X1 NOR2X1_1475 ( .A(_4201_), .B(_4198_), .Y(_4202_) );
NOR2X1 NOR2X1_1476 ( .A(_4202_), .B(_4200_), .Y(_0__26_) );
INVX1 INVX1_1379 ( .A(count_cycle_27_), .Y(_4203_) );
INVX1 INVX1_1380 ( .A(_4202_), .Y(_4204_) );
NOR2X1 NOR2X1_1477 ( .A(_4201_), .B(_4203_), .Y(_4205_) );
INVX1 INVX1_1381 ( .A(_4205_), .Y(_4206_) );
OAI21X1 OAI21X1_4301 ( .A(_4198_), .B(_4206_), .C(resetn_bF_buf10), .Y(_4207_) );
AOI21X1 AOI21X1_1068 ( .A(_4203_), .B(_4204_), .C(_4207_), .Y(_0__27_) );
NOR2X1 NOR2X1_1478 ( .A(_4196_), .B(_4206_), .Y(_4208_) );
NAND2X1 NAND2X1_1436 ( .A(_4208_), .B(_4189_), .Y(_4209_) );
INVX1 INVX1_1382 ( .A(_4209_), .Y(_4210_) );
OAI21X1 OAI21X1_4302 ( .A(_4210_), .B(count_cycle_28_), .C(resetn_bF_buf9), .Y(_4211_) );
INVX1 INVX1_1383 ( .A(count_cycle_28_), .Y(_4212_) );
NOR2X1 NOR2X1_1479 ( .A(_4212_), .B(_4209_), .Y(_4213_) );
NOR2X1 NOR2X1_1480 ( .A(_4213_), .B(_4211_), .Y(_0__28_) );
NOR2X1 NOR2X1_1481 ( .A(count_cycle_29_), .B(_4213_), .Y(_4214_) );
NAND2X1 NAND2X1_1437 ( .A(_4205_), .B(_4199_), .Y(_4215_) );
AND2X2 AND2X2_276 ( .A(count_cycle_28_), .B(count_cycle_29_), .Y(_4216_) );
INVX1 INVX1_1384 ( .A(_4216_), .Y(_4217_) );
OAI21X1 OAI21X1_4303 ( .A(_4215_), .B(_4217_), .C(resetn_bF_buf8), .Y(_4218_) );
NOR2X1 NOR2X1_1482 ( .A(_4214_), .B(_4218_), .Y(_0__29_) );
NOR2X1 NOR2X1_1483 ( .A(_4217_), .B(_4215_), .Y(_4219_) );
OAI21X1 OAI21X1_4304 ( .A(_4219_), .B(count_cycle_30_), .C(resetn_bF_buf7), .Y(_4220_) );
AOI21X1 AOI21X1_1069 ( .A(count_cycle_30_), .B(_4219_), .C(_4220_), .Y(_0__30_) );
AOI21X1 AOI21X1_1070 ( .A(count_cycle_30_), .B(_4219_), .C(count_cycle_31_), .Y(_4221_) );
OR2X2 OR2X2_52 ( .A(_4180_), .B(_4186_), .Y(_4222_) );
NOR2X1 NOR2X1_1484 ( .A(_4170_), .B(_4222_), .Y(_4223_) );
NAND2X1 NAND2X1_1438 ( .A(count_cycle_30_), .B(count_cycle_31_), .Y(_4224_) );
NOR2X1 NOR2X1_1485 ( .A(_4224_), .B(_4217_), .Y(_4225_) );
NAND3X1 NAND3X1_116 ( .A(_4208_), .B(_4225_), .C(_4223_), .Y(_4226_) );
OAI21X1 OAI21X1_4305 ( .A(_4163_), .B(_4226_), .C(resetn_bF_buf6), .Y(_4227_) );
NOR2X1 NOR2X1_1486 ( .A(_4227_), .B(_4221_), .Y(_0__31_) );
NOR2X1 NOR2X1_1487 ( .A(_4226_), .B(_4163_), .Y(_4228_) );
OAI21X1 OAI21X1_4306 ( .A(_4228_), .B(count_cycle_32_), .C(resetn_bF_buf5), .Y(_4229_) );
AOI21X1 AOI21X1_1071 ( .A(count_cycle_32_), .B(_4228_), .C(_4229_), .Y(_0__32_) );
INVX1 INVX1_1385 ( .A(count_cycle_33_), .Y(_4230_) );
NAND2X1 NAND2X1_1439 ( .A(count_cycle_32_), .B(_4228_), .Y(_4231_) );
OAI21X1 OAI21X1_4307 ( .A(_4231_), .B(_4230_), .C(resetn_bF_buf4), .Y(_4232_) );
AOI21X1 AOI21X1_1072 ( .A(_4230_), .B(_4231_), .C(_4232_), .Y(_0__33_) );
NOR2X1 NOR2X1_1488 ( .A(_4230_), .B(_4231_), .Y(_4233_) );
AND2X2 AND2X2_277 ( .A(_4233_), .B(count_cycle_34_), .Y(_4234_) );
OAI21X1 OAI21X1_4308 ( .A(_4233_), .B(count_cycle_34_), .C(resetn_bF_buf3), .Y(_4235_) );
NOR2X1 NOR2X1_1489 ( .A(_4235_), .B(_4234_), .Y(_0__34_) );
NAND2X1 NAND2X1_1440 ( .A(count_cycle_32_), .B(count_cycle_33_), .Y(_4236_) );
NAND2X1 NAND2X1_1441 ( .A(count_cycle_34_), .B(count_cycle_35_), .Y(_4237_) );
NOR2X1 NOR2X1_1490 ( .A(_4236_), .B(_4237_), .Y(_4238_) );
NAND2X1 NAND2X1_1442 ( .A(_4238_), .B(_4228_), .Y(_4239_) );
INVX1 INVX1_1386 ( .A(_4239_), .Y(_4240_) );
OAI21X1 OAI21X1_4309 ( .A(_4234_), .B(count_cycle_35_), .C(resetn_bF_buf2), .Y(_4241_) );
NOR2X1 NOR2X1_1491 ( .A(_4240_), .B(_4241_), .Y(_0__35_) );
INVX1 INVX1_1387 ( .A(count_cycle_36_), .Y(_4242_) );
NOR2X1 NOR2X1_1492 ( .A(_4242_), .B(_4239_), .Y(_4243_) );
OAI21X1 OAI21X1_4310 ( .A(_4240_), .B(count_cycle_36_), .C(resetn_bF_buf1), .Y(_4244_) );
NOR2X1 NOR2X1_1493 ( .A(_4243_), .B(_4244_), .Y(_0__36_) );
INVX1 INVX1_1388 ( .A(_4243_), .Y(_4245_) );
NOR2X1 NOR2X1_1494 ( .A(_4242_), .B(_2508_), .Y(_4246_) );
INVX1 INVX1_1389 ( .A(_4246_), .Y(_4247_) );
OAI21X1 OAI21X1_4311 ( .A(_4239_), .B(_4247_), .C(resetn_bF_buf0), .Y(_4248_) );
AOI21X1 AOI21X1_1073 ( .A(_2508_), .B(_4245_), .C(_4248_), .Y(_0__37_) );
NOR2X1 NOR2X1_1495 ( .A(_4247_), .B(_4239_), .Y(_4249_) );
OAI21X1 OAI21X1_4312 ( .A(_4249_), .B(count_cycle_38_), .C(resetn_bF_buf11), .Y(_4250_) );
AOI21X1 AOI21X1_1074 ( .A(count_cycle_38_), .B(_4249_), .C(_4250_), .Y(_0__38_) );
AOI21X1 AOI21X1_1075 ( .A(count_cycle_38_), .B(_4249_), .C(count_cycle_39_), .Y(_4251_) );
INVX1 INVX1_1390 ( .A(_4249_), .Y(_4252_) );
NAND2X1 NAND2X1_1443 ( .A(count_cycle_38_), .B(count_cycle_39_), .Y(_4253_) );
OAI21X1 OAI21X1_4313 ( .A(_4252_), .B(_4253_), .C(resetn_bF_buf10), .Y(_4254_) );
NOR2X1 NOR2X1_1496 ( .A(_4251_), .B(_4254_), .Y(_0__39_) );
NOR2X1 NOR2X1_1497 ( .A(_4253_), .B(_4247_), .Y(_4255_) );
AND2X2 AND2X2_278 ( .A(_4255_), .B(_4238_), .Y(_4256_) );
AND2X2 AND2X2_279 ( .A(_4228_), .B(_4256_), .Y(_4257_) );
OAI21X1 OAI21X1_4314 ( .A(_4257_), .B(count_cycle_40_), .C(resetn_bF_buf9), .Y(_4258_) );
AOI21X1 AOI21X1_1076 ( .A(count_cycle_40_), .B(_4257_), .C(_4258_), .Y(_0__40_) );
NAND2X1 NAND2X1_1444 ( .A(count_cycle_40_), .B(_4257_), .Y(_4259_) );
OAI21X1 OAI21X1_4315 ( .A(_4259_), .B(_2591_), .C(resetn_bF_buf8), .Y(_4260_) );
AOI21X1 AOI21X1_1077 ( .A(_2591_), .B(_4259_), .C(_4260_), .Y(_0__41_) );
NOR2X1 NOR2X1_1498 ( .A(_2591_), .B(_4259_), .Y(_4261_) );
AND2X2 AND2X2_280 ( .A(_4261_), .B(count_cycle_42_), .Y(_4262_) );
OAI21X1 OAI21X1_4316 ( .A(_4261_), .B(count_cycle_42_), .C(resetn_bF_buf7), .Y(_4263_) );
NOR2X1 NOR2X1_1499 ( .A(_4263_), .B(_4262_), .Y(_0__42_) );
NOR2X1 NOR2X1_1500 ( .A(count_cycle_43_), .B(_4262_), .Y(_4264_) );
NAND2X1 NAND2X1_1445 ( .A(count_cycle_40_), .B(count_cycle_41_), .Y(_4265_) );
NAND2X1 NAND2X1_1446 ( .A(count_cycle_42_), .B(count_cycle_43_), .Y(_4266_) );
NOR2X1 NOR2X1_1501 ( .A(_4265_), .B(_4266_), .Y(_4267_) );
NAND2X1 NAND2X1_1447 ( .A(_4267_), .B(_4257_), .Y(_4268_) );
NAND2X1 NAND2X1_1448 ( .A(resetn_bF_buf6), .B(_4268_), .Y(_4269_) );
NOR2X1 NOR2X1_1502 ( .A(_4269_), .B(_4264_), .Y(_0__43_) );
INVX1 INVX1_1391 ( .A(count_cycle_44_), .Y(_4270_) );
NOR2X1 NOR2X1_1503 ( .A(_4270_), .B(_4268_), .Y(_4271_) );
INVX1 INVX1_1392 ( .A(_4268_), .Y(_4272_) );
OAI21X1 OAI21X1_4317 ( .A(_4272_), .B(count_cycle_44_), .C(resetn_bF_buf5), .Y(_4273_) );
NOR2X1 NOR2X1_1504 ( .A(_4271_), .B(_4273_), .Y(_0__44_) );
INVX1 INVX1_1393 ( .A(count_cycle_45_), .Y(_4274_) );
OAI21X1 OAI21X1_4318 ( .A(_4268_), .B(_4270_), .C(_4274_), .Y(_4275_) );
NOR2X1 NOR2X1_1505 ( .A(_4270_), .B(_4274_), .Y(_4276_) );
INVX1 INVX1_1394 ( .A(_4276_), .Y(_4277_) );
OAI21X1 OAI21X1_4319 ( .A(_4268_), .B(_4277_), .C(_4275_), .Y(_4278_) );
NOR2X1 NOR2X1_1506 ( .A(_4426__bF_buf9), .B(_4278_), .Y(_0__45_) );
NAND3X1 NAND3X1_117 ( .A(count_cycle_46_), .B(_4276_), .C(_4272_), .Y(_4279_) );
OAI21X1 OAI21X1_4320 ( .A(_4268_), .B(_4277_), .C(_2691_), .Y(_4280_) );
AND2X2 AND2X2_281 ( .A(_4280_), .B(resetn_bF_buf4), .Y(_4281_) );
AND2X2 AND2X2_282 ( .A(_4281_), .B(_4279_), .Y(_0__46_) );
NAND2X1 NAND2X1_1449 ( .A(count_cycle_46_), .B(count_cycle_47_), .Y(_4282_) );
NOR2X1 NOR2X1_1507 ( .A(_4282_), .B(_4277_), .Y(_4283_) );
AND2X2 AND2X2_283 ( .A(_4283_), .B(_4267_), .Y(_4284_) );
AND2X2 AND2X2_284 ( .A(_4284_), .B(_4256_), .Y(_4285_) );
AND2X2 AND2X2_285 ( .A(_4228_), .B(_4285_), .Y(_4286_) );
INVX1 INVX1_1395 ( .A(_4286_), .Y(_4287_) );
NAND2X1 NAND2X1_1450 ( .A(resetn_bF_buf3), .B(_4287_), .Y(_4288_) );
AOI21X1 AOI21X1_1078 ( .A(_2706_), .B(_4279_), .C(_4288_), .Y(_0__47_) );
OAI21X1 OAI21X1_4321 ( .A(_4286_), .B(count_cycle_48_), .C(resetn_bF_buf2), .Y(_4289_) );
AOI21X1 AOI21X1_1079 ( .A(count_cycle_48_), .B(_4286_), .C(_4289_), .Y(_0__48_) );
INVX1 INVX1_1396 ( .A(count_cycle_48_), .Y(_4290_) );
OAI21X1 OAI21X1_4322 ( .A(_4287_), .B(_4290_), .C(_2756_), .Y(_4291_) );
NOR2X1 NOR2X1_1508 ( .A(_4290_), .B(_2756_), .Y(_4292_) );
INVX1 INVX1_1397 ( .A(_4292_), .Y(_4293_) );
OAI21X1 OAI21X1_4323 ( .A(_4287_), .B(_4293_), .C(_4291_), .Y(_4294_) );
NOR2X1 NOR2X1_1509 ( .A(_4426__bF_buf8), .B(_4294_), .Y(_0__49_) );
NOR2X1 NOR2X1_1510 ( .A(_4293_), .B(_4287_), .Y(_4295_) );
OAI21X1 OAI21X1_4324 ( .A(_4295_), .B(count_cycle_50_), .C(resetn_bF_buf1), .Y(_4296_) );
AOI21X1 AOI21X1_1080 ( .A(count_cycle_50_), .B(_4295_), .C(_4296_), .Y(_0__50_) );
NAND2X1 NAND2X1_1451 ( .A(count_cycle_50_), .B(_4295_), .Y(_4297_) );
NAND2X1 NAND2X1_1452 ( .A(count_cycle_50_), .B(count_cycle_51_), .Y(_4298_) );
NOR2X1 NOR2X1_1511 ( .A(_4298_), .B(_4293_), .Y(_4299_) );
NAND2X1 NAND2X1_1453 ( .A(_4299_), .B(_4286_), .Y(_4300_) );
NAND2X1 NAND2X1_1454 ( .A(resetn_bF_buf0), .B(_4300_), .Y(_4301_) );
AOI21X1 AOI21X1_1081 ( .A(_2786_), .B(_4297_), .C(_4301_), .Y(_0__51_) );
INVX1 INVX1_1398 ( .A(_4300_), .Y(_4302_) );
NAND2X1 NAND2X1_1455 ( .A(count_cycle_52_), .B(_4302_), .Y(_4303_) );
INVX1 INVX1_1399 ( .A(_4303_), .Y(_4304_) );
OAI21X1 OAI21X1_4325 ( .A(_4302_), .B(count_cycle_52_), .C(resetn_bF_buf11), .Y(_4305_) );
NOR2X1 NOR2X1_1512 ( .A(_4305_), .B(_4304_), .Y(_0__52_) );
INVX1 INVX1_1400 ( .A(count_cycle_53_), .Y(_4306_) );
NOR2X1 NOR2X1_1513 ( .A(_4306_), .B(_4303_), .Y(_4307_) );
OAI21X1 OAI21X1_4326 ( .A(_4304_), .B(count_cycle_53_), .C(resetn_bF_buf10), .Y(_4308_) );
NOR2X1 NOR2X1_1514 ( .A(_4307_), .B(_4308_), .Y(_0__53_) );
NAND2X1 NAND2X1_1456 ( .A(count_cycle_52_), .B(count_cycle_53_), .Y(_4309_) );
NOR2X1 NOR2X1_1515 ( .A(_4309_), .B(_4300_), .Y(_4310_) );
OAI21X1 OAI21X1_4327 ( .A(_4307_), .B(count_cycle_54_), .C(resetn_bF_buf9), .Y(_4311_) );
AOI21X1 AOI21X1_1082 ( .A(count_cycle_54_), .B(_4310_), .C(_4311_), .Y(_0__54_) );
AOI21X1 AOI21X1_1083 ( .A(count_cycle_54_), .B(_4310_), .C(count_cycle_55_), .Y(_4312_) );
NAND3X1 NAND3X1_118 ( .A(count_cycle_53_), .B(count_cycle_54_), .C(count_cycle_55_), .Y(_4313_) );
OAI21X1 OAI21X1_4328 ( .A(_4303_), .B(_4313_), .C(resetn_bF_buf8), .Y(_4314_) );
NOR2X1 NOR2X1_1516 ( .A(_4312_), .B(_4314_), .Y(_0__55_) );
NOR2X1 NOR2X1_1517 ( .A(_4313_), .B(_4303_), .Y(_4315_) );
OAI21X1 OAI21X1_4329 ( .A(_4315_), .B(count_cycle_56_), .C(resetn_bF_buf7), .Y(_4316_) );
AOI21X1 AOI21X1_1084 ( .A(count_cycle_56_), .B(_4315_), .C(_4316_), .Y(_0__56_) );
AOI21X1 AOI21X1_1085 ( .A(count_cycle_56_), .B(_4315_), .C(count_cycle_57_), .Y(_4317_) );
INVX1 INVX1_1401 ( .A(_4315_), .Y(_4318_) );
NAND2X1 NAND2X1_1457 ( .A(count_cycle_56_), .B(count_cycle_57_), .Y(_4319_) );
OAI21X1 OAI21X1_4330 ( .A(_4318_), .B(_4319_), .C(resetn_bF_buf6), .Y(_4320_) );
NOR2X1 NOR2X1_1518 ( .A(_4317_), .B(_4320_), .Y(_0__57_) );
NAND3X1 NAND3X1_119 ( .A(count_cycle_54_), .B(count_cycle_55_), .C(_4310_), .Y(_4321_) );
OAI21X1 OAI21X1_4331 ( .A(_4321_), .B(_4319_), .C(count_cycle_58_), .Y(_4322_) );
INVX1 INVX1_1402 ( .A(count_cycle_58_), .Y(_4323_) );
NOR2X1 NOR2X1_1519 ( .A(_4319_), .B(_4321_), .Y(_4324_) );
NAND2X1 NAND2X1_1458 ( .A(_4323_), .B(_4324_), .Y(_4325_) );
AOI21X1 AOI21X1_1086 ( .A(_4322_), .B(_4325_), .C(_4426__bF_buf7), .Y(_0__58_) );
NAND2X1 NAND2X1_1459 ( .A(count_cycle_58_), .B(_4324_), .Y(_4326_) );
NAND2X1 NAND2X1_1460 ( .A(count_cycle_59_), .B(_4326_), .Y(_4327_) );
OR2X2 OR2X2_53 ( .A(_4326_), .B(count_cycle_59_), .Y(_4328_) );
AOI21X1 AOI21X1_1087 ( .A(_4327_), .B(_4328_), .C(_4426__bF_buf6), .Y(_0__59_) );
INVX1 INVX1_1403 ( .A(_4319_), .Y(_4329_) );
NAND3X1 NAND3X1_120 ( .A(count_cycle_58_), .B(count_cycle_59_), .C(_4329_), .Y(_4330_) );
OAI21X1 OAI21X1_4332 ( .A(_4321_), .B(_4330_), .C(count_cycle_60_), .Y(_4331_) );
NOR2X1 NOR2X1_1520 ( .A(_4330_), .B(_4321_), .Y(_4332_) );
NAND2X1 NAND2X1_1461 ( .A(_2953_), .B(_4332_), .Y(_4333_) );
AOI21X1 AOI21X1_1088 ( .A(_4331_), .B(_4333_), .C(_4426__bF_buf5), .Y(_0__60_) );
NAND2X1 NAND2X1_1462 ( .A(count_cycle_60_), .B(_4332_), .Y(_4334_) );
NAND2X1 NAND2X1_1463 ( .A(count_cycle_61_), .B(_4334_), .Y(_4335_) );
OR2X2 OR2X2_54 ( .A(_4334_), .B(count_cycle_61_), .Y(_4336_) );
AOI21X1 AOI21X1_1089 ( .A(_4335_), .B(_4336_), .C(_4426__bF_buf4), .Y(_0__61_) );
NOR2X1 NOR2X1_1521 ( .A(_2953_), .B(_2967_), .Y(_4337_) );
NAND2X1 NAND2X1_1464 ( .A(_4337_), .B(_4332_), .Y(_4338_) );
NAND2X1 NAND2X1_1465 ( .A(count_cycle_62_), .B(_4338_), .Y(_4339_) );
AND2X2 AND2X2_286 ( .A(_4332_), .B(_4337_), .Y(_4340_) );
NAND2X1 NAND2X1_1466 ( .A(_2983_), .B(_4340_), .Y(_4341_) );
AOI21X1 AOI21X1_1090 ( .A(_4339_), .B(_4341_), .C(_4426__bF_buf3), .Y(_0__62_) );
OAI21X1 OAI21X1_4333 ( .A(_4338_), .B(_2983_), .C(count_cycle_63_), .Y(_4342_) );
INVX1 INVX1_1404 ( .A(count_cycle_63_), .Y(_4343_) );
NAND3X1 NAND3X1_121 ( .A(count_cycle_62_), .B(_4343_), .C(_4340_), .Y(_4344_) );
AOI21X1 AOI21X1_1091 ( .A(_4342_), .B(_4344_), .C(_4426__bF_buf2), .Y(_0__63_) );
NAND2X1 NAND2X1_1467 ( .A(_5273_), .B(_4638_), .Y(_4345_) );
OAI21X1 OAI21X1_4334 ( .A(_5359_), .B(_4638_), .C(_4345_), .Y(_1115_) );
MUX2X1 MUX2X1_298 ( .A(_4933__bF_buf4), .B(_5432_), .S(_4638_), .Y(_1116_) );
MUX2X1 MUX2X1_299 ( .A(_4940__bF_buf4), .B(_5501_), .S(_4638_), .Y(_1117_) );
MUX2X1 MUX2X1_300 ( .A(_4948__bF_buf4), .B(_5573_), .S(_4638_), .Y(_1118_) );
NAND2X1 NAND2X1_1468 ( .A(_4638_), .B(_5279_), .Y(_4346_) );
OAI21X1 OAI21X1_4335 ( .A(_5644_), .B(_4638_), .C(_4346_), .Y(_1119_) );
AND2X2 AND2X2_287 ( .A(resetn_bF_buf5), .B(cpu_state_0_), .Y(_86_) );
OAI21X1 OAI21X1_4336 ( .A(_4448_), .B(_4450_), .C(latched_is_lh), .Y(_4347_) );
AOI21X1 AOI21X1_1092 ( .A(_2568_), .B(_7631__bF_buf5), .C(_7629__bF_buf1), .Y(_4348_) );
OAI21X1 OAI21X1_4337 ( .A(instr_lh), .B(_7631__bF_buf4), .C(_4348_), .Y(_4349_) );
AOI21X1 AOI21X1_1093 ( .A(_4347_), .B(_4349_), .C(_4426__bF_buf1), .Y(_65_) );
OAI21X1 OAI21X1_4338 ( .A(_4448_), .B(_4450_), .C(latched_is_lu), .Y(_4350_) );
AOI21X1 AOI21X1_1094 ( .A(_2567_), .B(_7631__bF_buf3), .C(_7629__bF_buf0), .Y(_4351_) );
OAI21X1 OAI21X1_4339 ( .A(is_lbu_lhu_lw), .B(_7631__bF_buf2), .C(_4351_), .Y(_4352_) );
AOI21X1 AOI21X1_1095 ( .A(_4350_), .B(_4352_), .C(_4426__bF_buf0), .Y(_66_) );
NAND2X1 NAND2X1_1469 ( .A(_5847_), .B(_4556_), .Y(_4353_) );
NOR2X1 NOR2X1_1522 ( .A(_5261_), .B(_5251_), .Y(_4354_) );
AND2X2 AND2X2_288 ( .A(_5262_), .B(_5264_), .Y(_4355_) );
NAND3X1 NAND3X1_122 ( .A(is_beq_bne_blt_bge_bltu_bgeu), .B(_4355_), .C(_4354_), .Y(_4356_) );
NAND3X1 NAND3X1_123 ( .A(cpu_state_3_bF_buf4_), .B(_4353_), .C(_4356_), .Y(_4357_) );
AOI22X1 AOI22X1_167 ( .A(latched_branch), .B(_7625_), .C(_10099__bF_buf2), .D(instr_jal_bF_buf0), .Y(_4358_) );
AOI21X1 AOI21X1_1096 ( .A(_4358_), .B(_4357_), .C(_4426__bF_buf11), .Y(_63_) );
NOR2X1 NOR2X1_1523 ( .A(latched_stalu_bF_buf1), .B(_5737_), .Y(_4359_) );
OAI21X1 OAI21X1_4340 ( .A(_4431__bF_buf7), .B(cpu_state_3_bF_buf3_), .C(resetn_bF_buf4), .Y(_4360_) );
NOR2X1 NOR2X1_1524 ( .A(_4360_), .B(_4359_), .Y(_68_) );
OAI21X1 OAI21X1_4341 ( .A(_4533_), .B(latched_store), .C(cpu_state_2_bF_buf4_), .Y(_4361_) );
OAI21X1 OAI21X1_4342 ( .A(_4639__bF_buf3), .B(_4449_), .C(_4361_), .Y(_4362_) );
AOI21X1 AOI21X1_1097 ( .A(cpu_state_3_bF_buf2_), .B(_4356_), .C(_4362_), .Y(_4363_) );
NAND3X1 NAND3X1_124 ( .A(_4538__bF_buf1), .B(_4449_), .C(_7625_), .Y(_4364_) );
AOI21X1 AOI21X1_1098 ( .A(_4364_), .B(_4363_), .C(_4426__bF_buf10), .Y(_69_) );
INVX1 INVX1_1405 ( .A(_4472_), .Y(_4365_) );
OAI21X1 OAI21X1_4343 ( .A(_4435_), .B(_4455_), .C(_4365_), .Y(_74_) );
NAND3X1 NAND3X1_125 ( .A(_4476_), .B(_7627_), .C(_7628_), .Y(_4366_) );
OAI22X1 OAI22X1_312 ( .A(_4427_), .B(_4455_), .C(_4454_), .D(_4366_), .Y(_72_) );
OR2X2 OR2X2_55 ( .A(_5266_), .B(_4556_), .Y(_4367_) );
OAI21X1 OAI21X1_4344 ( .A(_4445_), .B(_4426__bF_buf9), .C(_4475_), .Y(_4368_) );
AOI21X1 AOI21X1_1099 ( .A(_4368_), .B(_7697__bF_buf3), .C(_4984_), .Y(_4369_) );
INVX1 INVX1_1406 ( .A(_4368_), .Y(_4370_) );
OAI21X1 OAI21X1_4345 ( .A(_4430_), .B(_4552_), .C(_4565_), .Y(_4371_) );
NOR2X1 NOR2X1_1525 ( .A(is_slli_srli_srai), .B(_4561_), .Y(_4372_) );
OAI21X1 OAI21X1_4346 ( .A(_4984_), .B(_4572_), .C(_4592_), .Y(_4373_) );
AOI21X1 AOI21X1_1100 ( .A(mem_do_prefetch_bF_buf5), .B(_4568_), .C(_4373_), .Y(_4374_) );
NAND3X1 NAND3X1_126 ( .A(_4552_), .B(_4565_), .C(_4372_), .Y(_4375_) );
OAI22X1 OAI22X1_313 ( .A(_4984_), .B(_4372_), .C(_4375_), .D(_4374_), .Y(_4376_) );
OAI21X1 OAI21X1_4347 ( .A(_4376_), .B(_4371_), .C(cpu_state_2_bF_buf3_), .Y(_4377_) );
AOI21X1 AOI21X1_1101 ( .A(mem_do_prefetch_bF_buf4), .B(_4597__bF_buf3), .C(_4607_), .Y(_4378_) );
AOI21X1 AOI21X1_1102 ( .A(_4378_), .B(_4377_), .C(_4370_), .Y(_4379_) );
OAI21X1 OAI21X1_4348 ( .A(_4379_), .B(_4369_), .C(_4456_), .Y(_4380_) );
OAI21X1 OAI21X1_4349 ( .A(_4367_), .B(_4603_), .C(_4380_), .Y(_73_) );
NAND2X1 NAND2X1_1470 ( .A(_1561_), .B(_1769_), .Y(_4381_) );
OAI21X1 OAI21X1_4350 ( .A(_4985__bF_buf0), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(resetn_bF_buf3), .Y(_4382_) );
AOI21X1 AOI21X1_1103 ( .A(_4985__bF_buf8), .B(_4381_), .C(_4382_), .Y(_52_) );
OAI21X1 OAI21X1_4351 ( .A(_4503_), .B(is_beq_bne_blt_bge_bltu_bgeu), .C(resetn_bF_buf2), .Y(_4383_) );
NOR2X1 NOR2X1_1526 ( .A(_1547__bF_buf2), .B(_4383_), .Y(_53_) );
OAI21X1 OAI21X1_4352 ( .A(_4605__bF_buf4), .B(decoder_pseudo_trigger_bF_buf2), .C(instr_and), .Y(_4384_) );
NAND2X1 NAND2X1_1471 ( .A(mem_rdata_q_12_), .B(mem_rdata_q_13_), .Y(_4385_) );
OR2X2 OR2X2_56 ( .A(_4385_), .B(_1575_), .Y(_4386_) );
NOR2X1 NOR2X1_1527 ( .A(_1746_), .B(_1568_), .Y(_4387_) );
INVX1 INVX1_1407 ( .A(_4387_), .Y(_4388_) );
OAI21X1 OAI21X1_4353 ( .A(_4388_), .B(_4386_), .C(_4384_), .Y(_4389_) );
AND2X2 AND2X2_289 ( .A(_4389_), .B(resetn_bF_buf1), .Y(_11_) );
NOR2X1 NOR2X1_1528 ( .A(_1575_), .B(_1712_), .Y(_4390_) );
AOI22X1 AOI22X1_168 ( .A(instr_or), .B(_1566__bF_buf2), .C(_4387_), .D(_4390_), .Y(_4391_) );
NOR2X1 NOR2X1_1529 ( .A(_4426__bF_buf8), .B(_4391_), .Y(_28_) );
OAI21X1 OAI21X1_4354 ( .A(_4605__bF_buf3), .B(decoder_pseudo_trigger_bF_buf1), .C(instr_sra), .Y(_4392_) );
INVX1 INVX1_1408 ( .A(_1745_), .Y(_4393_) );
NOR2X1 NOR2X1_1530 ( .A(_1553_), .B(_1760_), .Y(_4394_) );
NAND2X1 NAND2X1_1472 ( .A(_4393_), .B(_4394_), .Y(_4395_) );
AOI21X1 AOI21X1_1104 ( .A(_4392_), .B(_4395_), .C(_4426__bF_buf7), .Y(_42_) );
NAND2X1 NAND2X1_1473 ( .A(_1747_), .B(_4394_), .Y(_4396_) );
OAI21X1 OAI21X1_4355 ( .A(_4605__bF_buf2), .B(decoder_pseudo_trigger_bF_buf0), .C(instr_srl), .Y(_4397_) );
AOI21X1 AOI21X1_1105 ( .A(_4397_), .B(_4396_), .C(_4426__bF_buf6), .Y(_44_) );
OAI21X1 OAI21X1_4356 ( .A(_4605__bF_buf1), .B(decoder_pseudo_trigger_bF_buf3), .C(instr_xor), .Y(_4398_) );
OAI21X1 OAI21X1_4357 ( .A(_4388_), .B(_1763_), .C(_4398_), .Y(_4399_) );
AND2X2 AND2X2_290 ( .A(_4399_), .B(resetn_bF_buf0), .Y(_48_) );
NOR2X1 NOR2X1_1531 ( .A(mem_rdata_q_14_), .B(_4385_), .Y(_4400_) );
AOI22X1 AOI22X1_169 ( .A(instr_sltu), .B(_1566__bF_buf1), .C(_4387_), .D(_4400_), .Y(_4401_) );
NOR2X1 NOR2X1_1532 ( .A(_4426__bF_buf5), .B(_4401_), .Y(_41_) );
AOI22X1 AOI22X1_170 ( .A(instr_slt), .B(_1566__bF_buf0), .C(_4387_), .D(_1713_), .Y(_4402_) );
NOR2X1 NOR2X1_1533 ( .A(_4426__bF_buf4), .B(_4402_), .Y(_38_) );
AOI22X1 AOI22X1_171 ( .A(instr_sll), .B(_1566__bF_buf3), .C(_4387_), .D(_1750_), .Y(_4403_) );
NOR2X1 NOR2X1_1534 ( .A(_4426__bF_buf3), .B(_4403_), .Y(_36_) );
OAI21X1 OAI21X1_4358 ( .A(_4605__bF_buf0), .B(decoder_pseudo_trigger_bF_buf2), .C(instr_sub_bF_buf0), .Y(_4404_) );
NOR2X1 NOR2X1_1535 ( .A(_1553_), .B(_1758_), .Y(_4405_) );
NAND2X1 NAND2X1_1474 ( .A(_4405_), .B(_4393_), .Y(_4406_) );
AOI21X1 AOI21X1_1106 ( .A(_4404_), .B(_4406_), .C(_4426__bF_buf2), .Y(_46_) );
NAND2X1 NAND2X1_1475 ( .A(_4405_), .B(_1747_), .Y(_4407_) );
OAI21X1 OAI21X1_4359 ( .A(_4605__bF_buf5), .B(decoder_pseudo_trigger_bF_buf1), .C(instr_add), .Y(_4408_) );
AOI21X1 AOI21X1_1107 ( .A(_4408_), .B(_4407_), .C(_4426__bF_buf1), .Y(_9_) );
OAI21X1 OAI21X1_4360 ( .A(_4605__bF_buf4), .B(decoder_pseudo_trigger_bF_buf0), .C(instr_andi), .Y(_4409_) );
OAI21X1 OAI21X1_4361 ( .A(_1585_), .B(_4386_), .C(_4409_), .Y(_4410_) );
AND2X2 AND2X2_291 ( .A(_4410_), .B(resetn_bF_buf11), .Y(_12_) );
AOI22X1 AOI22X1_172 ( .A(instr_ori), .B(_1566__bF_buf2), .C(_1584_), .D(_4390_), .Y(_4411_) );
NOR2X1 NOR2X1_1536 ( .A(_4426__bF_buf0), .B(_4411_), .Y(_29_) );
OAI21X1 OAI21X1_4362 ( .A(_4605__bF_buf3), .B(decoder_pseudo_trigger_bF_buf3), .C(instr_xori), .Y(_4412_) );
OAI21X1 OAI21X1_4363 ( .A(_1585_), .B(_1763_), .C(_4412_), .Y(_4413_) );
AND2X2 AND2X2_292 ( .A(_4413_), .B(resetn_bF_buf10), .Y(_49_) );
AOI22X1 AOI22X1_173 ( .A(instr_sltiu), .B(_1566__bF_buf1), .C(_1584_), .D(_4400_), .Y(_4414_) );
NOR2X1 NOR2X1_1537 ( .A(_4426__bF_buf11), .B(_4414_), .Y(_40_) );
AOI22X1 AOI22X1_174 ( .A(instr_slti), .B(_1566__bF_buf0), .C(_1584_), .D(_1713_), .Y(_4415_) );
NOR2X1 NOR2X1_1538 ( .A(_4426__bF_buf10), .B(_4415_), .Y(_39_) );
AOI22X1 AOI22X1_175 ( .A(instr_addi), .B(_1566__bF_buf3), .C(_1584_), .D(_1757_), .Y(_4416_) );
NOR2X1 NOR2X1_1539 ( .A(_4426__bF_buf9), .B(_4416_), .Y(_10_) );
NOR2X1 NOR2X1_1540 ( .A(_4556_), .B(_1566__bF_buf2), .Y(_4417_) );
INVX1 INVX1_1409 ( .A(_4417_), .Y(_4418_) );
OAI22X1 OAI22X1_314 ( .A(_5252_), .B(_1547__bF_buf1), .C(_4418_), .D(_4386_), .Y(_4419_) );
AND2X2 AND2X2_293 ( .A(_4419_), .B(resetn_bF_buf9), .Y(_16_) );
AOI22X1 AOI22X1_176 ( .A(instr_bltu), .B(_1566__bF_buf1), .C(_4390_), .D(_4417_), .Y(_4420_) );
NOR2X1 NOR2X1_1541 ( .A(_4426__bF_buf8), .B(_4420_), .Y(_18_) );
AOI22X1 AOI22X1_177 ( .A(instr_bge), .B(_1566__bF_buf0), .C(_1742_), .D(_4417_), .Y(_4421_) );
NOR2X1 NOR2X1_1542 ( .A(_4426__bF_buf7), .B(_4421_), .Y(_15_) );
OAI22X1 OAI22X1_315 ( .A(_4522_), .B(_1547__bF_buf0), .C(_4418_), .D(_1763_), .Y(_4422_) );
AND2X2 AND2X2_294 ( .A(_4422_), .B(resetn_bF_buf8), .Y(_17_) );
AOI22X1 AOI22X1_178 ( .A(instr_bne), .B(_1566__bF_buf3), .C(_1750_), .D(_4417_), .Y(_4423_) );
NOR2X1 NOR2X1_1543 ( .A(_4426__bF_buf6), .B(_4423_), .Y(_19_) );
AOI22X1 AOI22X1_179 ( .A(instr_beq), .B(_1566__bF_buf2), .C(_4417_), .D(_1757_), .Y(_4424_) );
NOR2X1 NOR2X1_1544 ( .A(_4426__bF_buf5), .B(_4424_), .Y(_14_) );
BUFX2 BUFX2_1343 ( .A(cpuregs_0_[0]), .Y(_346_) );
BUFX2 BUFX2_1344 ( .A(cpuregs_0_[1]), .Y(_347_) );
BUFX2 BUFX2_1345 ( .A(cpuregs_0_[2]), .Y(_348_) );
BUFX2 BUFX2_1346 ( .A(cpuregs_0_[3]), .Y(_349_) );
BUFX2 BUFX2_1347 ( .A(cpuregs_0_[4]), .Y(_350_) );
BUFX2 BUFX2_1348 ( .A(cpuregs_0_[5]), .Y(_351_) );
BUFX2 BUFX2_1349 ( .A(cpuregs_0_[6]), .Y(_352_) );
BUFX2 BUFX2_1350 ( .A(cpuregs_0_[7]), .Y(_353_) );
BUFX2 BUFX2_1351 ( .A(cpuregs_0_[8]), .Y(_354_) );
BUFX2 BUFX2_1352 ( .A(cpuregs_0_[9]), .Y(_355_) );
BUFX2 BUFX2_1353 ( .A(cpuregs_0_[10]), .Y(_356_) );
BUFX2 BUFX2_1354 ( .A(cpuregs_0_[11]), .Y(_357_) );
BUFX2 BUFX2_1355 ( .A(cpuregs_0_[12]), .Y(_358_) );
BUFX2 BUFX2_1356 ( .A(cpuregs_0_[13]), .Y(_359_) );
BUFX2 BUFX2_1357 ( .A(cpuregs_0_[14]), .Y(_360_) );
BUFX2 BUFX2_1358 ( .A(cpuregs_0_[15]), .Y(_361_) );
BUFX2 BUFX2_1359 ( .A(cpuregs_0_[16]), .Y(_362_) );
BUFX2 BUFX2_1360 ( .A(cpuregs_0_[17]), .Y(_363_) );
BUFX2 BUFX2_1361 ( .A(cpuregs_0_[18]), .Y(_364_) );
BUFX2 BUFX2_1362 ( .A(cpuregs_0_[19]), .Y(_365_) );
BUFX2 BUFX2_1363 ( .A(cpuregs_0_[20]), .Y(_366_) );
BUFX2 BUFX2_1364 ( .A(cpuregs_0_[21]), .Y(_367_) );
BUFX2 BUFX2_1365 ( .A(cpuregs_0_[22]), .Y(_368_) );
BUFX2 BUFX2_1366 ( .A(cpuregs_0_[23]), .Y(_369_) );
BUFX2 BUFX2_1367 ( .A(cpuregs_0_[24]), .Y(_370_) );
BUFX2 BUFX2_1368 ( .A(cpuregs_0_[25]), .Y(_371_) );
BUFX2 BUFX2_1369 ( .A(cpuregs_0_[26]), .Y(_372_) );
BUFX2 BUFX2_1370 ( .A(cpuregs_0_[27]), .Y(_373_) );
BUFX2 BUFX2_1371 ( .A(cpuregs_0_[28]), .Y(_374_) );
BUFX2 BUFX2_1372 ( .A(cpuregs_0_[29]), .Y(_375_) );
BUFX2 BUFX2_1373 ( .A(cpuregs_0_[30]), .Y(_376_) );
BUFX2 BUFX2_1374 ( .A(cpuregs_0_[31]), .Y(_377_) );
BUFX2 BUFX2_1375 ( .A(gnd), .Y(eoi[0]) );
BUFX2 BUFX2_1376 ( .A(gnd), .Y(eoi[1]) );
BUFX2 BUFX2_1377 ( .A(gnd), .Y(eoi[2]) );
BUFX2 BUFX2_1378 ( .A(gnd), .Y(eoi[3]) );
BUFX2 BUFX2_1379 ( .A(gnd), .Y(eoi[4]) );
BUFX2 BUFX2_1380 ( .A(gnd), .Y(eoi[5]) );
BUFX2 BUFX2_1381 ( .A(gnd), .Y(eoi[6]) );
BUFX2 BUFX2_1382 ( .A(gnd), .Y(eoi[7]) );
BUFX2 BUFX2_1383 ( .A(gnd), .Y(eoi[8]) );
BUFX2 BUFX2_1384 ( .A(gnd), .Y(eoi[9]) );
BUFX2 BUFX2_1385 ( .A(gnd), .Y(eoi[10]) );
BUFX2 BUFX2_1386 ( .A(gnd), .Y(eoi[11]) );
BUFX2 BUFX2_1387 ( .A(gnd), .Y(eoi[12]) );
BUFX2 BUFX2_1388 ( .A(gnd), .Y(eoi[13]) );
BUFX2 BUFX2_1389 ( .A(gnd), .Y(eoi[14]) );
BUFX2 BUFX2_1390 ( .A(gnd), .Y(eoi[15]) );
BUFX2 BUFX2_1391 ( .A(gnd), .Y(eoi[16]) );
BUFX2 BUFX2_1392 ( .A(gnd), .Y(eoi[17]) );
BUFX2 BUFX2_1393 ( .A(gnd), .Y(eoi[18]) );
BUFX2 BUFX2_1394 ( .A(gnd), .Y(eoi[19]) );
BUFX2 BUFX2_1395 ( .A(gnd), .Y(eoi[20]) );
BUFX2 BUFX2_1396 ( .A(gnd), .Y(eoi[21]) );
BUFX2 BUFX2_1397 ( .A(gnd), .Y(eoi[22]) );
BUFX2 BUFX2_1398 ( .A(gnd), .Y(eoi[23]) );
BUFX2 BUFX2_1399 ( .A(gnd), .Y(eoi[24]) );
BUFX2 BUFX2_1400 ( .A(gnd), .Y(eoi[25]) );
BUFX2 BUFX2_1401 ( .A(gnd), .Y(eoi[26]) );
BUFX2 BUFX2_1402 ( .A(gnd), .Y(eoi[27]) );
BUFX2 BUFX2_1403 ( .A(gnd), .Y(eoi[28]) );
BUFX2 BUFX2_1404 ( .A(gnd), .Y(eoi[29]) );
BUFX2 BUFX2_1405 ( .A(gnd), .Y(eoi[30]) );
BUFX2 BUFX2_1406 ( .A(gnd), .Y(eoi[31]) );
BUFX2 BUFX2_1407 ( .A(_10724__0_), .Y(mem_addr[0]) );
BUFX2 BUFX2_1408 ( .A(_10724__1_), .Y(mem_addr[1]) );
BUFX2 BUFX2_1409 ( .A(_10724__2_), .Y(mem_addr[2]) );
BUFX2 BUFX2_1410 ( .A(_10724__3_), .Y(mem_addr[3]) );
BUFX2 BUFX2_1411 ( .A(_10724__4_), .Y(mem_addr[4]) );
BUFX2 BUFX2_1412 ( .A(_10724__5_), .Y(mem_addr[5]) );
BUFX2 BUFX2_1413 ( .A(_10724__6_), .Y(mem_addr[6]) );
BUFX2 BUFX2_1414 ( .A(_10724__7_), .Y(mem_addr[7]) );
BUFX2 BUFX2_1415 ( .A(_10724__8_), .Y(mem_addr[8]) );
BUFX2 BUFX2_1416 ( .A(_10724__9_), .Y(mem_addr[9]) );
BUFX2 BUFX2_1417 ( .A(_10724__10_), .Y(mem_addr[10]) );
BUFX2 BUFX2_1418 ( .A(_10724__11_), .Y(mem_addr[11]) );
BUFX2 BUFX2_1419 ( .A(_10724__12_), .Y(mem_addr[12]) );
BUFX2 BUFX2_1420 ( .A(_10724__13_), .Y(mem_addr[13]) );
BUFX2 BUFX2_1421 ( .A(_10724__14_), .Y(mem_addr[14]) );
BUFX2 BUFX2_1422 ( .A(_10724__15_), .Y(mem_addr[15]) );
BUFX2 BUFX2_1423 ( .A(_10724__16_), .Y(mem_addr[16]) );
BUFX2 BUFX2_1424 ( .A(_10724__17_), .Y(mem_addr[17]) );
BUFX2 BUFX2_1425 ( .A(_10724__18_), .Y(mem_addr[18]) );
BUFX2 BUFX2_1426 ( .A(_10724__19_), .Y(mem_addr[19]) );
BUFX2 BUFX2_1427 ( .A(_10724__20_), .Y(mem_addr[20]) );
BUFX2 BUFX2_1428 ( .A(_10724__21_), .Y(mem_addr[21]) );
BUFX2 BUFX2_1429 ( .A(_10724__22_), .Y(mem_addr[22]) );
BUFX2 BUFX2_1430 ( .A(_10724__23_), .Y(mem_addr[23]) );
BUFX2 BUFX2_1431 ( .A(_10724__24_), .Y(mem_addr[24]) );
BUFX2 BUFX2_1432 ( .A(_10724__25_), .Y(mem_addr[25]) );
BUFX2 BUFX2_1433 ( .A(_10724__26_), .Y(mem_addr[26]) );
BUFX2 BUFX2_1434 ( .A(_10724__27_), .Y(mem_addr[27]) );
BUFX2 BUFX2_1435 ( .A(_10724__28_), .Y(mem_addr[28]) );
BUFX2 BUFX2_1436 ( .A(_10724__29_), .Y(mem_addr[29]) );
BUFX2 BUFX2_1437 ( .A(_10724__30_), .Y(mem_addr[30]) );
BUFX2 BUFX2_1438 ( .A(_10724__31_), .Y(mem_addr[31]) );
BUFX2 BUFX2_1439 ( .A(_10725_), .Y(mem_instr) );
BUFX2 BUFX2_1440 ( .A(gnd), .Y(mem_la_addr[0]) );
BUFX2 BUFX2_1441 ( .A(gnd), .Y(mem_la_addr[1]) );
BUFX2 BUFX2_1442 ( .A(_10726__2_), .Y(mem_la_addr[2]) );
BUFX2 BUFX2_1443 ( .A(_10726__3_), .Y(mem_la_addr[3]) );
BUFX2 BUFX2_1444 ( .A(_10726__4_), .Y(mem_la_addr[4]) );
BUFX2 BUFX2_1445 ( .A(_10726__5_), .Y(mem_la_addr[5]) );
BUFX2 BUFX2_1446 ( .A(_10726__6_), .Y(mem_la_addr[6]) );
BUFX2 BUFX2_1447 ( .A(_10726__7_), .Y(mem_la_addr[7]) );
BUFX2 BUFX2_1448 ( .A(_10726__8_), .Y(mem_la_addr[8]) );
BUFX2 BUFX2_1449 ( .A(_10726__9_), .Y(mem_la_addr[9]) );
BUFX2 BUFX2_1450 ( .A(_10726__10_), .Y(mem_la_addr[10]) );
BUFX2 BUFX2_1451 ( .A(_10726__11_), .Y(mem_la_addr[11]) );
BUFX2 BUFX2_1452 ( .A(_10726__12_), .Y(mem_la_addr[12]) );
BUFX2 BUFX2_1453 ( .A(_10726__13_), .Y(mem_la_addr[13]) );
BUFX2 BUFX2_1454 ( .A(_10726__14_), .Y(mem_la_addr[14]) );
BUFX2 BUFX2_1455 ( .A(_10726__15_), .Y(mem_la_addr[15]) );
BUFX2 BUFX2_1456 ( .A(_10726__16_), .Y(mem_la_addr[16]) );
BUFX2 BUFX2_1457 ( .A(_10726__17_), .Y(mem_la_addr[17]) );
BUFX2 BUFX2_1458 ( .A(_10726__18_), .Y(mem_la_addr[18]) );
BUFX2 BUFX2_1459 ( .A(_10726__19_), .Y(mem_la_addr[19]) );
BUFX2 BUFX2_1460 ( .A(_10726__20_), .Y(mem_la_addr[20]) );
BUFX2 BUFX2_1461 ( .A(_10726__21_), .Y(mem_la_addr[21]) );
BUFX2 BUFX2_1462 ( .A(_10726__22_), .Y(mem_la_addr[22]) );
BUFX2 BUFX2_1463 ( .A(_10726__23_), .Y(mem_la_addr[23]) );
BUFX2 BUFX2_1464 ( .A(_10726__24_), .Y(mem_la_addr[24]) );
BUFX2 BUFX2_1465 ( .A(_10726__25_), .Y(mem_la_addr[25]) );
BUFX2 BUFX2_1466 ( .A(_10726__26_), .Y(mem_la_addr[26]) );
BUFX2 BUFX2_1467 ( .A(_10726__27_), .Y(mem_la_addr[27]) );
BUFX2 BUFX2_1468 ( .A(_10726__28_), .Y(mem_la_addr[28]) );
BUFX2 BUFX2_1469 ( .A(_10726__29_), .Y(mem_la_addr[29]) );
BUFX2 BUFX2_1470 ( .A(_10726__30_), .Y(mem_la_addr[30]) );
BUFX2 BUFX2_1471 ( .A(_10726__31_), .Y(mem_la_addr[31]) );
BUFX2 BUFX2_1472 ( .A(_10727_), .Y(mem_la_read) );
BUFX2 BUFX2_1473 ( .A(_10728__0_bF_buf4_), .Y(mem_la_wdata[0]) );
BUFX2 BUFX2_1474 ( .A(_10728__1_bF_buf0_), .Y(mem_la_wdata[1]) );
BUFX2 BUFX2_1475 ( .A(_10728__2_bF_buf4_), .Y(mem_la_wdata[2]) );
BUFX2 BUFX2_1476 ( .A(_10728__3_bF_buf3_), .Y(mem_la_wdata[3]) );
BUFX2 BUFX2_1477 ( .A(_10728__4_bF_buf0_), .Y(mem_la_wdata[4]) );
BUFX2 BUFX2_1478 ( .A(_10728__5_), .Y(mem_la_wdata[5]) );
BUFX2 BUFX2_1479 ( .A(_10728__6_), .Y(mem_la_wdata[6]) );
BUFX2 BUFX2_1480 ( .A(_10728__7_), .Y(mem_la_wdata[7]) );
BUFX2 BUFX2_1481 ( .A(_10728__8_), .Y(mem_la_wdata[8]) );
BUFX2 BUFX2_1482 ( .A(_10728__9_), .Y(mem_la_wdata[9]) );
BUFX2 BUFX2_1483 ( .A(_10728__10_), .Y(mem_la_wdata[10]) );
BUFX2 BUFX2_1484 ( .A(_10728__11_), .Y(mem_la_wdata[11]) );
BUFX2 BUFX2_1485 ( .A(_10728__12_), .Y(mem_la_wdata[12]) );
BUFX2 BUFX2_1486 ( .A(_10728__13_), .Y(mem_la_wdata[13]) );
BUFX2 BUFX2_1487 ( .A(_10728__14_), .Y(mem_la_wdata[14]) );
BUFX2 BUFX2_1488 ( .A(_10728__15_), .Y(mem_la_wdata[15]) );
BUFX2 BUFX2_1489 ( .A(_10728__16_), .Y(mem_la_wdata[16]) );
BUFX2 BUFX2_1490 ( .A(_10728__17_), .Y(mem_la_wdata[17]) );
BUFX2 BUFX2_1491 ( .A(_10728__18_), .Y(mem_la_wdata[18]) );
BUFX2 BUFX2_1492 ( .A(_10728__19_), .Y(mem_la_wdata[19]) );
BUFX2 BUFX2_1493 ( .A(_10728__20_), .Y(mem_la_wdata[20]) );
BUFX2 BUFX2_1494 ( .A(_10728__21_), .Y(mem_la_wdata[21]) );
BUFX2 BUFX2_1495 ( .A(_10728__22_), .Y(mem_la_wdata[22]) );
BUFX2 BUFX2_1496 ( .A(_10728__23_), .Y(mem_la_wdata[23]) );
BUFX2 BUFX2_1497 ( .A(_10728__24_), .Y(mem_la_wdata[24]) );
BUFX2 BUFX2_1498 ( .A(_10728__25_), .Y(mem_la_wdata[25]) );
BUFX2 BUFX2_1499 ( .A(_10728__26_), .Y(mem_la_wdata[26]) );
BUFX2 BUFX2_1500 ( .A(_10728__27_), .Y(mem_la_wdata[27]) );
BUFX2 BUFX2_1501 ( .A(_10728__28_), .Y(mem_la_wdata[28]) );
BUFX2 BUFX2_1502 ( .A(_10728__29_), .Y(mem_la_wdata[29]) );
BUFX2 BUFX2_1503 ( .A(_10728__30_), .Y(mem_la_wdata[30]) );
BUFX2 BUFX2_1504 ( .A(_10728__31_), .Y(mem_la_wdata[31]) );
BUFX2 BUFX2_1505 ( .A(_10729_), .Y(mem_la_write) );
BUFX2 BUFX2_1506 ( .A(_10730__0_), .Y(mem_la_wstrb[0]) );
BUFX2 BUFX2_1507 ( .A(_10730__1_), .Y(mem_la_wstrb[1]) );
BUFX2 BUFX2_1508 ( .A(_10730__2_), .Y(mem_la_wstrb[2]) );
BUFX2 BUFX2_1509 ( .A(_10730__3_), .Y(mem_la_wstrb[3]) );
BUFX2 BUFX2_1510 ( .A(_10731_), .Y(mem_valid) );
BUFX2 BUFX2_1511 ( .A(_10732__0_), .Y(mem_wdata[0]) );
BUFX2 BUFX2_1512 ( .A(_10732__1_), .Y(mem_wdata[1]) );
BUFX2 BUFX2_1513 ( .A(_10732__2_), .Y(mem_wdata[2]) );
BUFX2 BUFX2_1514 ( .A(_10732__3_), .Y(mem_wdata[3]) );
BUFX2 BUFX2_1515 ( .A(_10732__4_), .Y(mem_wdata[4]) );
BUFX2 BUFX2_1516 ( .A(_10732__5_), .Y(mem_wdata[5]) );
BUFX2 BUFX2_1517 ( .A(_10732__6_), .Y(mem_wdata[6]) );
BUFX2 BUFX2_1518 ( .A(_10732__7_), .Y(mem_wdata[7]) );
BUFX2 BUFX2_1519 ( .A(_10732__8_), .Y(mem_wdata[8]) );
BUFX2 BUFX2_1520 ( .A(_10732__9_), .Y(mem_wdata[9]) );
BUFX2 BUFX2_1521 ( .A(_10732__10_), .Y(mem_wdata[10]) );
BUFX2 BUFX2_1522 ( .A(_10732__11_), .Y(mem_wdata[11]) );
BUFX2 BUFX2_1523 ( .A(_10732__12_), .Y(mem_wdata[12]) );
BUFX2 BUFX2_1524 ( .A(_10732__13_), .Y(mem_wdata[13]) );
BUFX2 BUFX2_1525 ( .A(_10732__14_), .Y(mem_wdata[14]) );
BUFX2 BUFX2_1526 ( .A(_10732__15_), .Y(mem_wdata[15]) );
BUFX2 BUFX2_1527 ( .A(_10732__16_), .Y(mem_wdata[16]) );
BUFX2 BUFX2_1528 ( .A(_10732__17_), .Y(mem_wdata[17]) );
BUFX2 BUFX2_1529 ( .A(_10732__18_), .Y(mem_wdata[18]) );
BUFX2 BUFX2_1530 ( .A(_10732__19_), .Y(mem_wdata[19]) );
BUFX2 BUFX2_1531 ( .A(_10732__20_), .Y(mem_wdata[20]) );
BUFX2 BUFX2_1532 ( .A(_10732__21_), .Y(mem_wdata[21]) );
BUFX2 BUFX2_1533 ( .A(_10732__22_), .Y(mem_wdata[22]) );
BUFX2 BUFX2_1534 ( .A(_10732__23_), .Y(mem_wdata[23]) );
BUFX2 BUFX2_1535 ( .A(_10732__24_), .Y(mem_wdata[24]) );
BUFX2 BUFX2_1536 ( .A(_10732__25_), .Y(mem_wdata[25]) );
BUFX2 BUFX2_1537 ( .A(_10732__26_), .Y(mem_wdata[26]) );
BUFX2 BUFX2_1538 ( .A(_10732__27_), .Y(mem_wdata[27]) );
BUFX2 BUFX2_1539 ( .A(_10732__28_), .Y(mem_wdata[28]) );
BUFX2 BUFX2_1540 ( .A(_10732__29_), .Y(mem_wdata[29]) );
BUFX2 BUFX2_1541 ( .A(_10732__30_), .Y(mem_wdata[30]) );
BUFX2 BUFX2_1542 ( .A(_10732__31_), .Y(mem_wdata[31]) );
BUFX2 BUFX2_1543 ( .A(_10733__0_), .Y(mem_wstrb[0]) );
BUFX2 BUFX2_1544 ( .A(_10733__1_), .Y(mem_wstrb[1]) );
BUFX2 BUFX2_1545 ( .A(_10733__2_), .Y(mem_wstrb[2]) );
BUFX2 BUFX2_1546 ( .A(_10733__3_), .Y(mem_wstrb[3]) );
BUFX2 BUFX2_1547 ( .A(_undef), .Y(pcpi_insn[0]) );
BUFX2 BUFX2_1548 ( .A(_undef), .Y(pcpi_insn[1]) );
BUFX2 BUFX2_1549 ( .A(_undef), .Y(pcpi_insn[2]) );
BUFX2 BUFX2_1550 ( .A(_undef), .Y(pcpi_insn[3]) );
BUFX2 BUFX2_1551 ( .A(_undef), .Y(pcpi_insn[4]) );
BUFX2 BUFX2_1552 ( .A(_undef), .Y(pcpi_insn[5]) );
BUFX2 BUFX2_1553 ( .A(_undef), .Y(pcpi_insn[6]) );
BUFX2 BUFX2_1554 ( .A(_undef), .Y(pcpi_insn[7]) );
BUFX2 BUFX2_1555 ( .A(_undef), .Y(pcpi_insn[8]) );
BUFX2 BUFX2_1556 ( .A(_undef), .Y(pcpi_insn[9]) );
BUFX2 BUFX2_1557 ( .A(_undef), .Y(pcpi_insn[10]) );
BUFX2 BUFX2_1558 ( .A(_undef), .Y(pcpi_insn[11]) );
BUFX2 BUFX2_1559 ( .A(_undef), .Y(pcpi_insn[12]) );
BUFX2 BUFX2_1560 ( .A(_undef), .Y(pcpi_insn[13]) );
BUFX2 BUFX2_1561 ( .A(_undef), .Y(pcpi_insn[14]) );
BUFX2 BUFX2_1562 ( .A(_undef), .Y(pcpi_insn[15]) );
BUFX2 BUFX2_1563 ( .A(_undef), .Y(pcpi_insn[16]) );
BUFX2 BUFX2_1564 ( .A(_undef), .Y(pcpi_insn[17]) );
BUFX2 BUFX2_1565 ( .A(_undef), .Y(pcpi_insn[18]) );
BUFX2 BUFX2_1566 ( .A(_undef), .Y(pcpi_insn[19]) );
BUFX2 BUFX2_1567 ( .A(_undef), .Y(pcpi_insn[20]) );
BUFX2 BUFX2_1568 ( .A(_undef), .Y(pcpi_insn[21]) );
BUFX2 BUFX2_1569 ( .A(_undef), .Y(pcpi_insn[22]) );
BUFX2 BUFX2_1570 ( .A(_undef), .Y(pcpi_insn[23]) );
BUFX2 BUFX2_1571 ( .A(_undef), .Y(pcpi_insn[24]) );
BUFX2 BUFX2_1572 ( .A(_undef), .Y(pcpi_insn[25]) );
BUFX2 BUFX2_1573 ( .A(_undef), .Y(pcpi_insn[26]) );
BUFX2 BUFX2_1574 ( .A(_undef), .Y(pcpi_insn[27]) );
BUFX2 BUFX2_1575 ( .A(_undef), .Y(pcpi_insn[28]) );
BUFX2 BUFX2_1576 ( .A(_undef), .Y(pcpi_insn[29]) );
BUFX2 BUFX2_1577 ( .A(_undef), .Y(pcpi_insn[30]) );
BUFX2 BUFX2_1578 ( .A(_undef), .Y(pcpi_insn[31]) );
BUFX2 BUFX2_1579 ( .A(_10734__0_), .Y(pcpi_rs1[0]) );
BUFX2 BUFX2_1580 ( .A(_10734__1_), .Y(pcpi_rs1[1]) );
BUFX2 BUFX2_1581 ( .A(_10734__2_), .Y(pcpi_rs1[2]) );
BUFX2 BUFX2_1582 ( .A(_10734__3_), .Y(pcpi_rs1[3]) );
BUFX2 BUFX2_1583 ( .A(_10734__4_), .Y(pcpi_rs1[4]) );
BUFX2 BUFX2_1584 ( .A(_10734__5_), .Y(pcpi_rs1[5]) );
BUFX2 BUFX2_1585 ( .A(_10734__6_), .Y(pcpi_rs1[6]) );
BUFX2 BUFX2_1586 ( .A(_10734__7_), .Y(pcpi_rs1[7]) );
BUFX2 BUFX2_1587 ( .A(_10734__8_), .Y(pcpi_rs1[8]) );
BUFX2 BUFX2_1588 ( .A(_10734__9_), .Y(pcpi_rs1[9]) );
BUFX2 BUFX2_1589 ( .A(_10734__10_), .Y(pcpi_rs1[10]) );
BUFX2 BUFX2_1590 ( .A(_10734__11_), .Y(pcpi_rs1[11]) );
BUFX2 BUFX2_1591 ( .A(_10734__12_), .Y(pcpi_rs1[12]) );
BUFX2 BUFX2_1592 ( .A(_10734__13_), .Y(pcpi_rs1[13]) );
BUFX2 BUFX2_1593 ( .A(_10734__14_), .Y(pcpi_rs1[14]) );
BUFX2 BUFX2_1594 ( .A(_10734__15_), .Y(pcpi_rs1[15]) );
BUFX2 BUFX2_1595 ( .A(_10734__16_), .Y(pcpi_rs1[16]) );
BUFX2 BUFX2_1596 ( .A(_10734__17_), .Y(pcpi_rs1[17]) );
BUFX2 BUFX2_1597 ( .A(_10734__18_), .Y(pcpi_rs1[18]) );
BUFX2 BUFX2_1598 ( .A(_10734__19_), .Y(pcpi_rs1[19]) );
BUFX2 BUFX2_1599 ( .A(_10734__20_), .Y(pcpi_rs1[20]) );
BUFX2 BUFX2_1600 ( .A(_10734__21_), .Y(pcpi_rs1[21]) );
BUFX2 BUFX2_1601 ( .A(_10734__22_), .Y(pcpi_rs1[22]) );
BUFX2 BUFX2_1602 ( .A(_10734__23_), .Y(pcpi_rs1[23]) );
BUFX2 BUFX2_1603 ( .A(_10734__24_), .Y(pcpi_rs1[24]) );
BUFX2 BUFX2_1604 ( .A(_10734__25_), .Y(pcpi_rs1[25]) );
BUFX2 BUFX2_1605 ( .A(_10734__26_), .Y(pcpi_rs1[26]) );
BUFX2 BUFX2_1606 ( .A(_10734__27_), .Y(pcpi_rs1[27]) );
BUFX2 BUFX2_1607 ( .A(_10734__28_), .Y(pcpi_rs1[28]) );
BUFX2 BUFX2_1608 ( .A(_10734__29_), .Y(pcpi_rs1[29]) );
BUFX2 BUFX2_1609 ( .A(_10734__30_), .Y(pcpi_rs1[30]) );
BUFX2 BUFX2_1610 ( .A(_10734__31_), .Y(pcpi_rs1[31]) );
BUFX2 BUFX2_1611 ( .A(_10728__0_bF_buf3_), .Y(pcpi_rs2[0]) );
BUFX2 BUFX2_1612 ( .A(_10728__1_bF_buf3_), .Y(pcpi_rs2[1]) );
BUFX2 BUFX2_1613 ( .A(_10728__2_bF_buf3_), .Y(pcpi_rs2[2]) );
BUFX2 BUFX2_1614 ( .A(_10728__3_bF_buf2_), .Y(pcpi_rs2[3]) );
BUFX2 BUFX2_1615 ( .A(_10728__4_bF_buf4_), .Y(pcpi_rs2[4]) );
BUFX2 BUFX2_1616 ( .A(_10728__5_), .Y(pcpi_rs2[5]) );
BUFX2 BUFX2_1617 ( .A(_10728__6_), .Y(pcpi_rs2[6]) );
BUFX2 BUFX2_1618 ( .A(_10728__7_), .Y(pcpi_rs2[7]) );
BUFX2 BUFX2_1619 ( .A(_10735__8_), .Y(pcpi_rs2[8]) );
BUFX2 BUFX2_1620 ( .A(_10735__9_), .Y(pcpi_rs2[9]) );
BUFX2 BUFX2_1621 ( .A(_10735__10_), .Y(pcpi_rs2[10]) );
BUFX2 BUFX2_1622 ( .A(_10735__11_), .Y(pcpi_rs2[11]) );
BUFX2 BUFX2_1623 ( .A(_10735__12_), .Y(pcpi_rs2[12]) );
BUFX2 BUFX2_1624 ( .A(_10735__13_), .Y(pcpi_rs2[13]) );
BUFX2 BUFX2_1625 ( .A(_10735__14_), .Y(pcpi_rs2[14]) );
BUFX2 BUFX2_1626 ( .A(_10735__15_), .Y(pcpi_rs2[15]) );
BUFX2 BUFX2_1627 ( .A(_10735__16_), .Y(pcpi_rs2[16]) );
BUFX2 BUFX2_1628 ( .A(_10735__17_), .Y(pcpi_rs2[17]) );
BUFX2 BUFX2_1629 ( .A(_10735__18_), .Y(pcpi_rs2[18]) );
BUFX2 BUFX2_1630 ( .A(_10735__19_), .Y(pcpi_rs2[19]) );
BUFX2 BUFX2_1631 ( .A(_10735__20_), .Y(pcpi_rs2[20]) );
BUFX2 BUFX2_1632 ( .A(_10735__21_), .Y(pcpi_rs2[21]) );
BUFX2 BUFX2_1633 ( .A(_10735__22_), .Y(pcpi_rs2[22]) );
BUFX2 BUFX2_1634 ( .A(_10735__23_), .Y(pcpi_rs2[23]) );
BUFX2 BUFX2_1635 ( .A(_10735__24_), .Y(pcpi_rs2[24]) );
BUFX2 BUFX2_1636 ( .A(_10735__25_), .Y(pcpi_rs2[25]) );
BUFX2 BUFX2_1637 ( .A(_10735__26_), .Y(pcpi_rs2[26]) );
BUFX2 BUFX2_1638 ( .A(_10735__27_), .Y(pcpi_rs2[27]) );
BUFX2 BUFX2_1639 ( .A(_10735__28_), .Y(pcpi_rs2[28]) );
BUFX2 BUFX2_1640 ( .A(_10735__29_), .Y(pcpi_rs2[29]) );
BUFX2 BUFX2_1641 ( .A(_10735__30_), .Y(pcpi_rs2[30]) );
BUFX2 BUFX2_1642 ( .A(_10735__31_), .Y(pcpi_rs2[31]) );
BUFX2 BUFX2_1643 ( .A(gnd), .Y(pcpi_valid) );
BUFX2 BUFX2_1644 ( .A(_undef), .Y(trace_data[0]) );
BUFX2 BUFX2_1645 ( .A(_undef), .Y(trace_data[1]) );
BUFX2 BUFX2_1646 ( .A(_undef), .Y(trace_data[2]) );
BUFX2 BUFX2_1647 ( .A(_undef), .Y(trace_data[3]) );
BUFX2 BUFX2_1648 ( .A(_undef), .Y(trace_data[4]) );
BUFX2 BUFX2_1649 ( .A(_undef), .Y(trace_data[5]) );
BUFX2 BUFX2_1650 ( .A(_undef), .Y(trace_data[6]) );
BUFX2 BUFX2_1651 ( .A(_undef), .Y(trace_data[7]) );
BUFX2 BUFX2_1652 ( .A(_undef), .Y(trace_data[8]) );
BUFX2 BUFX2_1653 ( .A(_undef), .Y(trace_data[9]) );
BUFX2 BUFX2_1654 ( .A(_undef), .Y(trace_data[10]) );
BUFX2 BUFX2_1655 ( .A(_undef), .Y(trace_data[11]) );
BUFX2 BUFX2_1656 ( .A(_undef), .Y(trace_data[12]) );
BUFX2 BUFX2_1657 ( .A(_undef), .Y(trace_data[13]) );
BUFX2 BUFX2_1658 ( .A(_undef), .Y(trace_data[14]) );
BUFX2 BUFX2_1659 ( .A(_undef), .Y(trace_data[15]) );
BUFX2 BUFX2_1660 ( .A(_undef), .Y(trace_data[16]) );
BUFX2 BUFX2_1661 ( .A(_undef), .Y(trace_data[17]) );
BUFX2 BUFX2_1662 ( .A(_undef), .Y(trace_data[18]) );
BUFX2 BUFX2_1663 ( .A(_undef), .Y(trace_data[19]) );
BUFX2 BUFX2_1664 ( .A(_undef), .Y(trace_data[20]) );
BUFX2 BUFX2_1665 ( .A(_undef), .Y(trace_data[21]) );
BUFX2 BUFX2_1666 ( .A(_undef), .Y(trace_data[22]) );
BUFX2 BUFX2_1667 ( .A(_undef), .Y(trace_data[23]) );
BUFX2 BUFX2_1668 ( .A(_undef), .Y(trace_data[24]) );
BUFX2 BUFX2_1669 ( .A(_undef), .Y(trace_data[25]) );
BUFX2 BUFX2_1670 ( .A(_undef), .Y(trace_data[26]) );
BUFX2 BUFX2_1671 ( .A(_undef), .Y(trace_data[27]) );
BUFX2 BUFX2_1672 ( .A(_undef), .Y(trace_data[28]) );
BUFX2 BUFX2_1673 ( .A(_undef), .Y(trace_data[29]) );
BUFX2 BUFX2_1674 ( .A(_undef), .Y(trace_data[30]) );
BUFX2 BUFX2_1675 ( .A(_undef), .Y(trace_data[31]) );
BUFX2 BUFX2_1676 ( .A(gnd), .Y(trace_data[32]) );
BUFX2 BUFX2_1677 ( .A(gnd), .Y(trace_data[33]) );
BUFX2 BUFX2_1678 ( .A(gnd), .Y(trace_data[34]) );
BUFX2 BUFX2_1679 ( .A(gnd), .Y(trace_data[35]) );
BUFX2 BUFX2_1680 ( .A(gnd), .Y(trace_valid) );
BUFX2 BUFX2_1681 ( .A(_10736_), .Y(trap) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf136), .D(_218_), .Q(cpuregs_4_[0]) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf135), .D(_219_), .Q(cpuregs_4_[1]) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf134), .D(_220_), .Q(cpuregs_4_[2]) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf133), .D(_221_), .Q(cpuregs_4_[3]) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf132), .D(_222_), .Q(cpuregs_4_[4]) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf131), .D(_223_), .Q(cpuregs_4_[5]) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf130), .D(_224_), .Q(cpuregs_4_[6]) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf129), .D(_225_), .Q(cpuregs_4_[7]) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf128), .D(_226_), .Q(cpuregs_4_[8]) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf127), .D(_227_), .Q(cpuregs_4_[9]) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf126), .D(_228_), .Q(cpuregs_4_[10]) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf125), .D(_229_), .Q(cpuregs_4_[11]) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf124), .D(_230_), .Q(cpuregs_4_[12]) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf123), .D(_231_), .Q(cpuregs_4_[13]) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf122), .D(_232_), .Q(cpuregs_4_[14]) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf121), .D(_233_), .Q(cpuregs_4_[15]) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf120), .D(_234_), .Q(cpuregs_4_[16]) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf119), .D(_235_), .Q(cpuregs_4_[17]) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf118), .D(_236_), .Q(cpuregs_4_[18]) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf117), .D(_237_), .Q(cpuregs_4_[19]) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf116), .D(_238_), .Q(cpuregs_4_[20]) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf115), .D(_239_), .Q(cpuregs_4_[21]) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf114), .D(_240_), .Q(cpuregs_4_[22]) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf113), .D(_241_), .Q(cpuregs_4_[23]) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf112), .D(_242_), .Q(cpuregs_4_[24]) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf111), .D(_243_), .Q(cpuregs_4_[25]) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf110), .D(_244_), .Q(cpuregs_4_[26]) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf109), .D(_245_), .Q(cpuregs_4_[27]) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf108), .D(_246_), .Q(cpuregs_4_[28]) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf107), .D(_247_), .Q(cpuregs_4_[29]) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf106), .D(_248_), .Q(cpuregs_4_[30]) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf105), .D(_249_), .Q(cpuregs_4_[31]) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf104), .D(_859_), .Q(cpuregs_19_[0]) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf103), .D(_860_), .Q(cpuregs_19_[1]) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf102), .D(_861_), .Q(cpuregs_19_[2]) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf101), .D(_862_), .Q(cpuregs_19_[3]) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf100), .D(_863_), .Q(cpuregs_19_[4]) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf99), .D(_864_), .Q(cpuregs_19_[5]) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf98), .D(_865_), .Q(cpuregs_19_[6]) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf97), .D(_866_), .Q(cpuregs_19_[7]) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf96), .D(_867_), .Q(cpuregs_19_[8]) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf95), .D(_868_), .Q(cpuregs_19_[9]) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf94), .D(_869_), .Q(cpuregs_19_[10]) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf93), .D(_870_), .Q(cpuregs_19_[11]) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf92), .D(_871_), .Q(cpuregs_19_[12]) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf91), .D(_872_), .Q(cpuregs_19_[13]) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf90), .D(_873_), .Q(cpuregs_19_[14]) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf89), .D(_874_), .Q(cpuregs_19_[15]) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf88), .D(_875_), .Q(cpuregs_19_[16]) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf87), .D(_876_), .Q(cpuregs_19_[17]) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf86), .D(_877_), .Q(cpuregs_19_[18]) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf85), .D(_878_), .Q(cpuregs_19_[19]) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf84), .D(_879_), .Q(cpuregs_19_[20]) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf83), .D(_880_), .Q(cpuregs_19_[21]) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf82), .D(_881_), .Q(cpuregs_19_[22]) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf81), .D(_882_), .Q(cpuregs_19_[23]) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf80), .D(_883_), .Q(cpuregs_19_[24]) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf79), .D(_884_), .Q(cpuregs_19_[25]) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf78), .D(_885_), .Q(cpuregs_19_[26]) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf77), .D(_886_), .Q(cpuregs_19_[27]) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf76), .D(_887_), .Q(cpuregs_19_[28]) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf75), .D(_888_), .Q(cpuregs_19_[29]) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf74), .D(_889_), .Q(cpuregs_19_[30]) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf73), .D(_890_), .Q(cpuregs_19_[31]) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf72), .D(_635_), .Q(cpuregs_23_[0]) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf71), .D(_636_), .Q(cpuregs_23_[1]) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf70), .D(_637_), .Q(cpuregs_23_[2]) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf69), .D(_638_), .Q(cpuregs_23_[3]) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf68), .D(_639_), .Q(cpuregs_23_[4]) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf67), .D(_640_), .Q(cpuregs_23_[5]) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf66), .D(_641_), .Q(cpuregs_23_[6]) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf65), .D(_642_), .Q(cpuregs_23_[7]) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf64), .D(_643_), .Q(cpuregs_23_[8]) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf63), .D(_644_), .Q(cpuregs_23_[9]) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf62), .D(_645_), .Q(cpuregs_23_[10]) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf61), .D(_646_), .Q(cpuregs_23_[11]) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf60), .D(_647_), .Q(cpuregs_23_[12]) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf59), .D(_648_), .Q(cpuregs_23_[13]) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf58), .D(_649_), .Q(cpuregs_23_[14]) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf57), .D(_650_), .Q(cpuregs_23_[15]) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf56), .D(_651_), .Q(cpuregs_23_[16]) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf55), .D(_652_), .Q(cpuregs_23_[17]) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf54), .D(_653_), .Q(cpuregs_23_[18]) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf53), .D(_654_), .Q(cpuregs_23_[19]) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf52), .D(_655_), .Q(cpuregs_23_[20]) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf51), .D(_656_), .Q(cpuregs_23_[21]) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf50), .D(_657_), .Q(cpuregs_23_[22]) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf49), .D(_658_), .Q(cpuregs_23_[23]) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf48), .D(_659_), .Q(cpuregs_23_[24]) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf47), .D(_660_), .Q(cpuregs_23_[25]) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf46), .D(_661_), .Q(cpuregs_23_[26]) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf45), .D(_662_), .Q(cpuregs_23_[27]) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf44), .D(_663_), .Q(cpuregs_23_[28]) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf43), .D(_664_), .Q(cpuregs_23_[29]) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf42), .D(_665_), .Q(cpuregs_23_[30]) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf41), .D(_666_), .Q(cpuregs_23_[31]) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf40), .D(_603_), .Q(cpuregs_24_[0]) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf39), .D(_604_), .Q(cpuregs_24_[1]) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf38), .D(_605_), .Q(cpuregs_24_[2]) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf37), .D(_606_), .Q(cpuregs_24_[3]) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf36), .D(_607_), .Q(cpuregs_24_[4]) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf35), .D(_608_), .Q(cpuregs_24_[5]) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf34), .D(_609_), .Q(cpuregs_24_[6]) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf33), .D(_610_), .Q(cpuregs_24_[7]) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf32), .D(_611_), .Q(cpuregs_24_[8]) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf31), .D(_612_), .Q(cpuregs_24_[9]) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf30), .D(_613_), .Q(cpuregs_24_[10]) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf29), .D(_614_), .Q(cpuregs_24_[11]) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf28), .D(_615_), .Q(cpuregs_24_[12]) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf27), .D(_616_), .Q(cpuregs_24_[13]) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf26), .D(_617_), .Q(cpuregs_24_[14]) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf25), .D(_618_), .Q(cpuregs_24_[15]) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf24), .D(_619_), .Q(cpuregs_24_[16]) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf23), .D(_620_), .Q(cpuregs_24_[17]) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf22), .D(_621_), .Q(cpuregs_24_[18]) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf21), .D(_622_), .Q(cpuregs_24_[19]) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf20), .D(_623_), .Q(cpuregs_24_[20]) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf19), .D(_624_), .Q(cpuregs_24_[21]) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf18), .D(_625_), .Q(cpuregs_24_[22]) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf17), .D(_626_), .Q(cpuregs_24_[23]) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf16), .D(_627_), .Q(cpuregs_24_[24]) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf15), .D(_628_), .Q(cpuregs_24_[25]) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf14), .D(_629_), .Q(cpuregs_24_[26]) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf13), .D(_630_), .Q(cpuregs_24_[27]) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf12), .D(_631_), .Q(cpuregs_24_[28]) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf11), .D(_632_), .Q(cpuregs_24_[29]) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf10), .D(_633_), .Q(cpuregs_24_[30]) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf9), .D(_634_), .Q(cpuregs_24_[31]) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf8), .D(_891_), .Q(cpuregs_12_[0]) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf7), .D(_892_), .Q(cpuregs_12_[1]) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf6), .D(_893_), .Q(cpuregs_12_[2]) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf5), .D(_894_), .Q(cpuregs_12_[3]) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf4), .D(_895_), .Q(cpuregs_12_[4]) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf3), .D(_896_), .Q(cpuregs_12_[5]) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf2), .D(_897_), .Q(cpuregs_12_[6]) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf1), .D(_898_), .Q(cpuregs_12_[7]) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf0), .D(_899_), .Q(cpuregs_12_[8]) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf136), .D(_900_), .Q(cpuregs_12_[9]) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf135), .D(_901_), .Q(cpuregs_12_[10]) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf134), .D(_902_), .Q(cpuregs_12_[11]) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf133), .D(_903_), .Q(cpuregs_12_[12]) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf132), .D(_904_), .Q(cpuregs_12_[13]) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf131), .D(_905_), .Q(cpuregs_12_[14]) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf130), .D(_906_), .Q(cpuregs_12_[15]) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf129), .D(_907_), .Q(cpuregs_12_[16]) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf128), .D(_908_), .Q(cpuregs_12_[17]) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf127), .D(_909_), .Q(cpuregs_12_[18]) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf126), .D(_910_), .Q(cpuregs_12_[19]) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf125), .D(_911_), .Q(cpuregs_12_[20]) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf124), .D(_912_), .Q(cpuregs_12_[21]) );
DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf123), .D(_913_), .Q(cpuregs_12_[22]) );
DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf122), .D(_914_), .Q(cpuregs_12_[23]) );
DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf121), .D(_915_), .Q(cpuregs_12_[24]) );
DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf120), .D(_916_), .Q(cpuregs_12_[25]) );
DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf119), .D(_917_), .Q(cpuregs_12_[26]) );
DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf118), .D(_918_), .Q(cpuregs_12_[27]) );
DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf117), .D(_919_), .Q(cpuregs_12_[28]) );
DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf116), .D(_920_), .Q(cpuregs_12_[29]) );
DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf115), .D(_921_), .Q(cpuregs_12_[30]) );
DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf114), .D(_922_), .Q(cpuregs_12_[31]) );
DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf113), .D(_571_), .Q(cpuregs_25_[0]) );
DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf112), .D(_572_), .Q(cpuregs_25_[1]) );
DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf111), .D(_573_), .Q(cpuregs_25_[2]) );
DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf110), .D(_574_), .Q(cpuregs_25_[3]) );
DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf109), .D(_575_), .Q(cpuregs_25_[4]) );
DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf108), .D(_576_), .Q(cpuregs_25_[5]) );
DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf107), .D(_577_), .Q(cpuregs_25_[6]) );
DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf106), .D(_578_), .Q(cpuregs_25_[7]) );
DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf105), .D(_579_), .Q(cpuregs_25_[8]) );
DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf104), .D(_580_), .Q(cpuregs_25_[9]) );
DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf103), .D(_581_), .Q(cpuregs_25_[10]) );
DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf102), .D(_582_), .Q(cpuregs_25_[11]) );
DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf101), .D(_583_), .Q(cpuregs_25_[12]) );
DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf100), .D(_584_), .Q(cpuregs_25_[13]) );
DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf99), .D(_585_), .Q(cpuregs_25_[14]) );
DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf98), .D(_586_), .Q(cpuregs_25_[15]) );
DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf97), .D(_587_), .Q(cpuregs_25_[16]) );
DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf96), .D(_588_), .Q(cpuregs_25_[17]) );
DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf95), .D(_589_), .Q(cpuregs_25_[18]) );
DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf94), .D(_590_), .Q(cpuregs_25_[19]) );
DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf93), .D(_591_), .Q(cpuregs_25_[20]) );
DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf92), .D(_592_), .Q(cpuregs_25_[21]) );
DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf91), .D(_593_), .Q(cpuregs_25_[22]) );
DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf90), .D(_594_), .Q(cpuregs_25_[23]) );
DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf89), .D(_595_), .Q(cpuregs_25_[24]) );
DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf88), .D(_596_), .Q(cpuregs_25_[25]) );
DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf87), .D(_597_), .Q(cpuregs_25_[26]) );
DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf86), .D(_598_), .Q(cpuregs_25_[27]) );
DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf85), .D(_599_), .Q(cpuregs_25_[28]) );
DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf84), .D(_600_), .Q(cpuregs_25_[29]) );
DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf83), .D(_601_), .Q(cpuregs_25_[30]) );
DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf82), .D(_602_), .Q(cpuregs_25_[31]) );
DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf81), .D(_795_), .Q(cpuregs_11_[0]) );
DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf80), .D(_796_), .Q(cpuregs_11_[1]) );
DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf79), .D(_797_), .Q(cpuregs_11_[2]) );
DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf78), .D(_798_), .Q(cpuregs_11_[3]) );
DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf77), .D(_799_), .Q(cpuregs_11_[4]) );
DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf76), .D(_800_), .Q(cpuregs_11_[5]) );
DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf75), .D(_801_), .Q(cpuregs_11_[6]) );
DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf74), .D(_802_), .Q(cpuregs_11_[7]) );
DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf73), .D(_803_), .Q(cpuregs_11_[8]) );
DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf72), .D(_804_), .Q(cpuregs_11_[9]) );
DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf71), .D(_805_), .Q(cpuregs_11_[10]) );
DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf70), .D(_806_), .Q(cpuregs_11_[11]) );
DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf69), .D(_807_), .Q(cpuregs_11_[12]) );
DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf68), .D(_808_), .Q(cpuregs_11_[13]) );
DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf67), .D(_809_), .Q(cpuregs_11_[14]) );
DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf66), .D(_810_), .Q(cpuregs_11_[15]) );
DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf65), .D(_811_), .Q(cpuregs_11_[16]) );
DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf64), .D(_812_), .Q(cpuregs_11_[17]) );
DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf63), .D(_813_), .Q(cpuregs_11_[18]) );
DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf62), .D(_814_), .Q(cpuregs_11_[19]) );
DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf61), .D(_815_), .Q(cpuregs_11_[20]) );
DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf60), .D(_816_), .Q(cpuregs_11_[21]) );
DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf59), .D(_817_), .Q(cpuregs_11_[22]) );
DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf58), .D(_818_), .Q(cpuregs_11_[23]) );
DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf57), .D(_819_), .Q(cpuregs_11_[24]) );
DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf56), .D(_820_), .Q(cpuregs_11_[25]) );
DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf55), .D(_821_), .Q(cpuregs_11_[26]) );
DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf54), .D(_822_), .Q(cpuregs_11_[27]) );
DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf53), .D(_823_), .Q(cpuregs_11_[28]) );
DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf52), .D(_824_), .Q(cpuregs_11_[29]) );
DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf51), .D(_825_), .Q(cpuregs_11_[30]) );
DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf50), .D(_826_), .Q(cpuregs_11_[31]) );
DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf49), .D(_763_), .Q(cpuregs_9_[0]) );
DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf48), .D(_764_), .Q(cpuregs_9_[1]) );
DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf47), .D(_765_), .Q(cpuregs_9_[2]) );
DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf46), .D(_766_), .Q(cpuregs_9_[3]) );
DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf45), .D(_767_), .Q(cpuregs_9_[4]) );
DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf44), .D(_768_), .Q(cpuregs_9_[5]) );
DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf43), .D(_769_), .Q(cpuregs_9_[6]) );
DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf42), .D(_770_), .Q(cpuregs_9_[7]) );
DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf41), .D(_771_), .Q(cpuregs_9_[8]) );
DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf40), .D(_772_), .Q(cpuregs_9_[9]) );
DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf39), .D(_773_), .Q(cpuregs_9_[10]) );
DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf38), .D(_774_), .Q(cpuregs_9_[11]) );
DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf37), .D(_775_), .Q(cpuregs_9_[12]) );
DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf36), .D(_776_), .Q(cpuregs_9_[13]) );
DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf35), .D(_777_), .Q(cpuregs_9_[14]) );
DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf34), .D(_778_), .Q(cpuregs_9_[15]) );
DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf33), .D(_779_), .Q(cpuregs_9_[16]) );
DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf32), .D(_780_), .Q(cpuregs_9_[17]) );
DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf31), .D(_781_), .Q(cpuregs_9_[18]) );
DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf30), .D(_782_), .Q(cpuregs_9_[19]) );
DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf29), .D(_783_), .Q(cpuregs_9_[20]) );
DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf28), .D(_784_), .Q(cpuregs_9_[21]) );
DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf27), .D(_785_), .Q(cpuregs_9_[22]) );
DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf26), .D(_786_), .Q(cpuregs_9_[23]) );
DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf25), .D(_787_), .Q(cpuregs_9_[24]) );
DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf24), .D(_788_), .Q(cpuregs_9_[25]) );
DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf23), .D(_789_), .Q(cpuregs_9_[26]) );
DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf22), .D(_790_), .Q(cpuregs_9_[27]) );
DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf21), .D(_791_), .Q(cpuregs_9_[28]) );
DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf20), .D(_792_), .Q(cpuregs_9_[29]) );
DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf19), .D(_793_), .Q(cpuregs_9_[30]) );
DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf18), .D(_794_), .Q(cpuregs_9_[31]) );
DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf17), .D(_539_), .Q(cpuregs_26_[0]) );
DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf16), .D(_540_), .Q(cpuregs_26_[1]) );
DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf15), .D(_541_), .Q(cpuregs_26_[2]) );
DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf14), .D(_542_), .Q(cpuregs_26_[3]) );
DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf13), .D(_543_), .Q(cpuregs_26_[4]) );
DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf12), .D(_544_), .Q(cpuregs_26_[5]) );
DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf11), .D(_545_), .Q(cpuregs_26_[6]) );
DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf10), .D(_546_), .Q(cpuregs_26_[7]) );
DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf9), .D(_547_), .Q(cpuregs_26_[8]) );
DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf8), .D(_548_), .Q(cpuregs_26_[9]) );
DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf7), .D(_549_), .Q(cpuregs_26_[10]) );
DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf6), .D(_550_), .Q(cpuregs_26_[11]) );
DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf5), .D(_551_), .Q(cpuregs_26_[12]) );
DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf4), .D(_552_), .Q(cpuregs_26_[13]) );
DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf3), .D(_553_), .Q(cpuregs_26_[14]) );
DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf2), .D(_554_), .Q(cpuregs_26_[15]) );
DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf1), .D(_555_), .Q(cpuregs_26_[16]) );
DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf0), .D(_556_), .Q(cpuregs_26_[17]) );
DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf136), .D(_557_), .Q(cpuregs_26_[18]) );
DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf135), .D(_558_), .Q(cpuregs_26_[19]) );
DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf134), .D(_559_), .Q(cpuregs_26_[20]) );
DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf133), .D(_560_), .Q(cpuregs_26_[21]) );
DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf132), .D(_561_), .Q(cpuregs_26_[22]) );
DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf131), .D(_562_), .Q(cpuregs_26_[23]) );
DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf130), .D(_563_), .Q(cpuregs_26_[24]) );
DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf129), .D(_564_), .Q(cpuregs_26_[25]) );
DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf128), .D(_565_), .Q(cpuregs_26_[26]) );
DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf127), .D(_566_), .Q(cpuregs_26_[27]) );
DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf126), .D(_567_), .Q(cpuregs_26_[28]) );
DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf125), .D(_568_), .Q(cpuregs_26_[29]) );
DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf124), .D(_569_), .Q(cpuregs_26_[30]) );
DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf123), .D(_570_), .Q(cpuregs_26_[31]) );
DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf122), .D(_411_), .Q(cpuregs_30_[0]) );
DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf121), .D(_412_), .Q(cpuregs_30_[1]) );
DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf120), .D(_413_), .Q(cpuregs_30_[2]) );
DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf119), .D(_414_), .Q(cpuregs_30_[3]) );
DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf118), .D(_415_), .Q(cpuregs_30_[4]) );
DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf117), .D(_416_), .Q(cpuregs_30_[5]) );
DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf116), .D(_417_), .Q(cpuregs_30_[6]) );
DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf115), .D(_418_), .Q(cpuregs_30_[7]) );
DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf114), .D(_419_), .Q(cpuregs_30_[8]) );
DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf113), .D(_420_), .Q(cpuregs_30_[9]) );
DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf112), .D(_421_), .Q(cpuregs_30_[10]) );
DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf111), .D(_422_), .Q(cpuregs_30_[11]) );
DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf110), .D(_423_), .Q(cpuregs_30_[12]) );
DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf109), .D(_424_), .Q(cpuregs_30_[13]) );
DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf108), .D(_425_), .Q(cpuregs_30_[14]) );
DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf107), .D(_426_), .Q(cpuregs_30_[15]) );
DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf106), .D(_427_), .Q(cpuregs_30_[16]) );
DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf105), .D(_428_), .Q(cpuregs_30_[17]) );
DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf104), .D(_429_), .Q(cpuregs_30_[18]) );
DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf103), .D(_430_), .Q(cpuregs_30_[19]) );
DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf102), .D(_431_), .Q(cpuregs_30_[20]) );
DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf101), .D(_432_), .Q(cpuregs_30_[21]) );
DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf100), .D(_433_), .Q(cpuregs_30_[22]) );
DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf99), .D(_434_), .Q(cpuregs_30_[23]) );
DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf98), .D(_435_), .Q(cpuregs_30_[24]) );
DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf97), .D(_436_), .Q(cpuregs_30_[25]) );
DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf96), .D(_437_), .Q(cpuregs_30_[26]) );
DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf95), .D(_438_), .Q(cpuregs_30_[27]) );
DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf94), .D(_439_), .Q(cpuregs_30_[28]) );
DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf93), .D(_440_), .Q(cpuregs_30_[29]) );
DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf92), .D(_441_), .Q(cpuregs_30_[30]) );
DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf91), .D(_442_), .Q(cpuregs_30_[31]) );
DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf90), .D(_379_), .Q(cpuregs_31_[0]) );
DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf89), .D(_380_), .Q(cpuregs_31_[1]) );
DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf88), .D(_381_), .Q(cpuregs_31_[2]) );
DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf87), .D(_382_), .Q(cpuregs_31_[3]) );
DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf86), .D(_383_), .Q(cpuregs_31_[4]) );
DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf85), .D(_384_), .Q(cpuregs_31_[5]) );
DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf84), .D(_385_), .Q(cpuregs_31_[6]) );
DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf83), .D(_386_), .Q(cpuregs_31_[7]) );
DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf82), .D(_387_), .Q(cpuregs_31_[8]) );
DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf81), .D(_388_), .Q(cpuregs_31_[9]) );
DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf80), .D(_389_), .Q(cpuregs_31_[10]) );
DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf79), .D(_390_), .Q(cpuregs_31_[11]) );
DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf78), .D(_391_), .Q(cpuregs_31_[12]) );
DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf77), .D(_392_), .Q(cpuregs_31_[13]) );
DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf76), .D(_393_), .Q(cpuregs_31_[14]) );
DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf75), .D(_394_), .Q(cpuregs_31_[15]) );
DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf74), .D(_395_), .Q(cpuregs_31_[16]) );
DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf73), .D(_396_), .Q(cpuregs_31_[17]) );
DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf72), .D(_397_), .Q(cpuregs_31_[18]) );
DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf71), .D(_398_), .Q(cpuregs_31_[19]) );
DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf70), .D(_399_), .Q(cpuregs_31_[20]) );
DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf69), .D(_400_), .Q(cpuregs_31_[21]) );
DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf68), .D(_401_), .Q(cpuregs_31_[22]) );
DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf67), .D(_402_), .Q(cpuregs_31_[23]) );
DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf66), .D(_403_), .Q(cpuregs_31_[24]) );
DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf65), .D(_404_), .Q(cpuregs_31_[25]) );
DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf64), .D(_405_), .Q(cpuregs_31_[26]) );
DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf63), .D(_406_), .Q(cpuregs_31_[27]) );
DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf62), .D(_407_), .Q(cpuregs_31_[28]) );
DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf61), .D(_408_), .Q(cpuregs_31_[29]) );
DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf60), .D(_409_), .Q(cpuregs_31_[30]) );
DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf59), .D(_410_), .Q(cpuregs_31_[31]) );
DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf58), .D(_5__0_), .Q(decoded_rs1_0_) );
DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf57), .D(_5__1_), .Q(decoded_rs1_1_) );
DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf56), .D(_5__2_), .Q(decoded_rs1_2_) );
DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf55), .D(_5__3_), .Q(decoded_rs1_3_) );
DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf54), .D(_5__4_), .Q(decoded_rs1_4_) );
DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf53), .D(_186_), .Q(cpuregs_5_[0]) );
DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf52), .D(_187_), .Q(cpuregs_5_[1]) );
DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf51), .D(_188_), .Q(cpuregs_5_[2]) );
DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf50), .D(_189_), .Q(cpuregs_5_[3]) );
DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf49), .D(_190_), .Q(cpuregs_5_[4]) );
DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf48), .D(_191_), .Q(cpuregs_5_[5]) );
DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf47), .D(_192_), .Q(cpuregs_5_[6]) );
DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf46), .D(_193_), .Q(cpuregs_5_[7]) );
DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf45), .D(_194_), .Q(cpuregs_5_[8]) );
DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf44), .D(_195_), .Q(cpuregs_5_[9]) );
DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf43), .D(_196_), .Q(cpuregs_5_[10]) );
DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf42), .D(_197_), .Q(cpuregs_5_[11]) );
DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf41), .D(_198_), .Q(cpuregs_5_[12]) );
DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf40), .D(_199_), .Q(cpuregs_5_[13]) );
DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf39), .D(_200_), .Q(cpuregs_5_[14]) );
DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf38), .D(_201_), .Q(cpuregs_5_[15]) );
DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf37), .D(_202_), .Q(cpuregs_5_[16]) );
DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf36), .D(_203_), .Q(cpuregs_5_[17]) );
DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf35), .D(_204_), .Q(cpuregs_5_[18]) );
DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf34), .D(_205_), .Q(cpuregs_5_[19]) );
DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf33), .D(_206_), .Q(cpuregs_5_[20]) );
DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf32), .D(_207_), .Q(cpuregs_5_[21]) );
DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf31), .D(_208_), .Q(cpuregs_5_[22]) );
DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf30), .D(_209_), .Q(cpuregs_5_[23]) );
DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf29), .D(_210_), .Q(cpuregs_5_[24]) );
DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf28), .D(_211_), .Q(cpuregs_5_[25]) );
DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf27), .D(_212_), .Q(cpuregs_5_[26]) );
DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf26), .D(_213_), .Q(cpuregs_5_[27]) );
DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf25), .D(_214_), .Q(cpuregs_5_[28]) );
DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf24), .D(_215_), .Q(cpuregs_5_[29]) );
DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf23), .D(_216_), .Q(cpuregs_5_[30]) );
DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf22), .D(_217_), .Q(cpuregs_5_[31]) );
DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf21), .D(_154_), .Q(cpuregs_6_[0]) );
DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf20), .D(_155_), .Q(cpuregs_6_[1]) );
DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf19), .D(_156_), .Q(cpuregs_6_[2]) );
DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf18), .D(_157_), .Q(cpuregs_6_[3]) );
DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf17), .D(_158_), .Q(cpuregs_6_[4]) );
DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf16), .D(_159_), .Q(cpuregs_6_[5]) );
DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf15), .D(_160_), .Q(cpuregs_6_[6]) );
DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf14), .D(_161_), .Q(cpuregs_6_[7]) );
DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf13), .D(_162_), .Q(cpuregs_6_[8]) );
DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf12), .D(_163_), .Q(cpuregs_6_[9]) );
DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf11), .D(_164_), .Q(cpuregs_6_[10]) );
DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf10), .D(_165_), .Q(cpuregs_6_[11]) );
DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf9), .D(_166_), .Q(cpuregs_6_[12]) );
DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf8), .D(_167_), .Q(cpuregs_6_[13]) );
DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf7), .D(_168_), .Q(cpuregs_6_[14]) );
DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf6), .D(_169_), .Q(cpuregs_6_[15]) );
DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf5), .D(_170_), .Q(cpuregs_6_[16]) );
DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf4), .D(_171_), .Q(cpuregs_6_[17]) );
DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf3), .D(_172_), .Q(cpuregs_6_[18]) );
DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf2), .D(_173_), .Q(cpuregs_6_[19]) );
DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf1), .D(_174_), .Q(cpuregs_6_[20]) );
DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf0), .D(_175_), .Q(cpuregs_6_[21]) );
DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf136), .D(_176_), .Q(cpuregs_6_[22]) );
DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf135), .D(_177_), .Q(cpuregs_6_[23]) );
DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf134), .D(_178_), .Q(cpuregs_6_[24]) );
DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf133), .D(_179_), .Q(cpuregs_6_[25]) );
DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf132), .D(_180_), .Q(cpuregs_6_[26]) );
DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf131), .D(_181_), .Q(cpuregs_6_[27]) );
DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf130), .D(_182_), .Q(cpuregs_6_[28]) );
DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf129), .D(_183_), .Q(cpuregs_6_[29]) );
DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf128), .D(_184_), .Q(cpuregs_6_[30]) );
DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf127), .D(_185_), .Q(cpuregs_6_[31]) );
DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf126), .D(_86_), .Q(_10736_) );
DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf125), .D(_0__0_), .Q(count_cycle_0_) );
DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf124), .D(_0__1_), .Q(count_cycle_1_) );
DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf123), .D(_0__2_), .Q(count_cycle_2_) );
DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf122), .D(_0__3_), .Q(count_cycle_3_) );
DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf121), .D(_0__4_), .Q(count_cycle_4_) );
DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf120), .D(_0__5_), .Q(count_cycle_5_) );
DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf119), .D(_0__6_), .Q(count_cycle_6_) );
DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf118), .D(_0__7_), .Q(count_cycle_7_) );
DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf117), .D(_0__8_), .Q(count_cycle_8_) );
DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf116), .D(_0__9_), .Q(count_cycle_9_) );
DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf115), .D(_0__10_), .Q(count_cycle_10_) );
DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf114), .D(_0__11_), .Q(count_cycle_11_) );
DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf113), .D(_0__12_), .Q(count_cycle_12_) );
DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf112), .D(_0__13_), .Q(count_cycle_13_) );
DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf111), .D(_0__14_), .Q(count_cycle_14_) );
DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf110), .D(_0__15_), .Q(count_cycle_15_) );
DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf109), .D(_0__16_), .Q(count_cycle_16_) );
DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf108), .D(_0__17_), .Q(count_cycle_17_) );
DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf107), .D(_0__18_), .Q(count_cycle_18_) );
DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf106), .D(_0__19_), .Q(count_cycle_19_) );
DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf105), .D(_0__20_), .Q(count_cycle_20_) );
DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf104), .D(_0__21_), .Q(count_cycle_21_) );
DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf103), .D(_0__22_), .Q(count_cycle_22_) );
DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf102), .D(_0__23_), .Q(count_cycle_23_) );
DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf101), .D(_0__24_), .Q(count_cycle_24_) );
DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf100), .D(_0__25_), .Q(count_cycle_25_) );
DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf99), .D(_0__26_), .Q(count_cycle_26_) );
DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf98), .D(_0__27_), .Q(count_cycle_27_) );
DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf97), .D(_0__28_), .Q(count_cycle_28_) );
DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf96), .D(_0__29_), .Q(count_cycle_29_) );
DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf95), .D(_0__30_), .Q(count_cycle_30_) );
DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf94), .D(_0__31_), .Q(count_cycle_31_) );
DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf93), .D(_0__32_), .Q(count_cycle_32_) );
DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf92), .D(_0__33_), .Q(count_cycle_33_) );
DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf91), .D(_0__34_), .Q(count_cycle_34_) );
DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf90), .D(_0__35_), .Q(count_cycle_35_) );
DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf89), .D(_0__36_), .Q(count_cycle_36_) );
DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf88), .D(_0__37_), .Q(count_cycle_37_) );
DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf87), .D(_0__38_), .Q(count_cycle_38_) );
DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf86), .D(_0__39_), .Q(count_cycle_39_) );
DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf85), .D(_0__40_), .Q(count_cycle_40_) );
DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf84), .D(_0__41_), .Q(count_cycle_41_) );
DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf83), .D(_0__42_), .Q(count_cycle_42_) );
DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf82), .D(_0__43_), .Q(count_cycle_43_) );
DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf81), .D(_0__44_), .Q(count_cycle_44_) );
DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf80), .D(_0__45_), .Q(count_cycle_45_) );
DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf79), .D(_0__46_), .Q(count_cycle_46_) );
DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf78), .D(_0__47_), .Q(count_cycle_47_) );
DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf77), .D(_0__48_), .Q(count_cycle_48_) );
DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf76), .D(_0__49_), .Q(count_cycle_49_) );
DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf75), .D(_0__50_), .Q(count_cycle_50_) );
DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf74), .D(_0__51_), .Q(count_cycle_51_) );
DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf73), .D(_0__52_), .Q(count_cycle_52_) );
DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf72), .D(_0__53_), .Q(count_cycle_53_) );
DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf71), .D(_0__54_), .Q(count_cycle_54_) );
DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf70), .D(_0__55_), .Q(count_cycle_55_) );
DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf69), .D(_0__56_), .Q(count_cycle_56_) );
DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf68), .D(_0__57_), .Q(count_cycle_57_) );
DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf67), .D(_0__58_), .Q(count_cycle_58_) );
DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf66), .D(_0__59_), .Q(count_cycle_59_) );
DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf65), .D(_0__60_), .Q(count_cycle_60_) );
DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf64), .D(_0__61_), .Q(count_cycle_61_) );
DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf63), .D(_0__62_), .Q(count_cycle_62_) );
DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf62), .D(_0__63_), .Q(count_cycle_63_) );
DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf61), .D(_1__0_), .Q(count_instr_0_) );
DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf60), .D(_1__1_), .Q(count_instr_1_) );
DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf59), .D(_1__2_), .Q(count_instr_2_) );
DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf58), .D(_1__3_), .Q(count_instr_3_) );
DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf57), .D(_1__4_), .Q(count_instr_4_) );
DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf56), .D(_1__5_), .Q(count_instr_5_) );
DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf55), .D(_1__6_), .Q(count_instr_6_) );
DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf54), .D(_1__7_), .Q(count_instr_7_) );
DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf53), .D(_1__8_), .Q(count_instr_8_) );
DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf52), .D(_1__9_), .Q(count_instr_9_) );
DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf51), .D(_1__10_), .Q(count_instr_10_) );
DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf50), .D(_1__11_), .Q(count_instr_11_) );
DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf49), .D(_1__12_), .Q(count_instr_12_) );
DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf48), .D(_1__13_), .Q(count_instr_13_) );
DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf47), .D(_1__14_), .Q(count_instr_14_) );
DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf46), .D(_1__15_), .Q(count_instr_15_) );
DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf45), .D(_1__16_), .Q(count_instr_16_) );
DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf44), .D(_1__17_), .Q(count_instr_17_) );
DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf43), .D(_1__18_), .Q(count_instr_18_) );
DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf42), .D(_1__19_), .Q(count_instr_19_) );
DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf41), .D(_1__20_), .Q(count_instr_20_) );
DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf40), .D(_1__21_), .Q(count_instr_21_) );
DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf39), .D(_1__22_), .Q(count_instr_22_) );
DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf38), .D(_1__23_), .Q(count_instr_23_) );
DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf37), .D(_1__24_), .Q(count_instr_24_) );
DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf36), .D(_1__25_), .Q(count_instr_25_) );
DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf35), .D(_1__26_), .Q(count_instr_26_) );
DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf34), .D(_1__27_), .Q(count_instr_27_) );
DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf33), .D(_1__28_), .Q(count_instr_28_) );
DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf32), .D(_1__29_), .Q(count_instr_29_) );
DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf31), .D(_1__30_), .Q(count_instr_30_) );
DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf30), .D(_1__31_), .Q(count_instr_31_) );
DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf29), .D(_1__32_), .Q(count_instr_32_) );
DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf28), .D(_1__33_), .Q(count_instr_33_) );
DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf27), .D(_1__34_), .Q(count_instr_34_) );
DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf26), .D(_1__35_), .Q(count_instr_35_) );
DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf25), .D(_1__36_), .Q(count_instr_36_) );
DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf24), .D(_1__37_), .Q(count_instr_37_) );
DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf23), .D(_1__38_), .Q(count_instr_38_) );
DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf22), .D(_1__39_), .Q(count_instr_39_) );
DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf21), .D(_1__40_), .Q(count_instr_40_) );
DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf20), .D(_1__41_), .Q(count_instr_41_) );
DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf19), .D(_1__42_), .Q(count_instr_42_) );
DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf18), .D(_1__43_), .Q(count_instr_43_) );
DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf17), .D(_1__44_), .Q(count_instr_44_) );
DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf16), .D(_1__45_), .Q(count_instr_45_) );
DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf15), .D(_1__46_), .Q(count_instr_46_) );
DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf14), .D(_1__47_), .Q(count_instr_47_) );
DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf13), .D(_1__48_), .Q(count_instr_48_) );
DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf12), .D(_1__49_), .Q(count_instr_49_) );
DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf11), .D(_1__50_), .Q(count_instr_50_) );
DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf10), .D(_1__51_), .Q(count_instr_51_) );
DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf9), .D(_1__52_), .Q(count_instr_52_) );
DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf8), .D(_1__53_), .Q(count_instr_53_) );
DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf7), .D(_1__54_), .Q(count_instr_54_) );
DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf6), .D(_1__55_), .Q(count_instr_55_) );
DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf5), .D(_1__56_), .Q(count_instr_56_) );
DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf4), .D(_1__57_), .Q(count_instr_57_) );
DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf3), .D(_1__58_), .Q(count_instr_58_) );
DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf2), .D(_1__59_), .Q(count_instr_59_) );
DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf1), .D(_1__60_), .Q(count_instr_60_) );
DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf0), .D(_1__61_), .Q(count_instr_61_) );
DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf136), .D(_1__62_), .Q(count_instr_62_) );
DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf135), .D(_1__63_), .Q(count_instr_63_) );
DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf134), .D(_84__0_), .Q(reg_pc_0_) );
DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf133), .D(_84__1_), .Q(reg_pc_1_) );
DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf132), .D(_84__2_), .Q(reg_pc_2_) );
DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf131), .D(_84__3_), .Q(reg_pc_3_) );
DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf130), .D(_84__4_), .Q(reg_pc_4_) );
DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf129), .D(_84__5_), .Q(reg_pc_5_) );
DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf128), .D(_84__6_), .Q(reg_pc_6_) );
DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf127), .D(_84__7_), .Q(reg_pc_7_) );
DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf126), .D(_84__8_), .Q(reg_pc_8_) );
DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf125), .D(_84__9_), .Q(reg_pc_9_) );
DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf124), .D(_84__10_), .Q(reg_pc_10_) );
DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf123), .D(_84__11_), .Q(reg_pc_11_) );
DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf122), .D(_84__12_), .Q(reg_pc_12_) );
DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf121), .D(_84__13_), .Q(reg_pc_13_) );
DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf120), .D(_84__14_), .Q(reg_pc_14_) );
DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf119), .D(_84__15_), .Q(reg_pc_15_) );
DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf118), .D(_84__16_), .Q(reg_pc_16_) );
DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf117), .D(_84__17_), .Q(reg_pc_17_) );
DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf116), .D(_84__18_), .Q(reg_pc_18_) );
DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf115), .D(_84__19_), .Q(reg_pc_19_) );
DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf114), .D(_84__20_), .Q(reg_pc_20_) );
DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf113), .D(_84__21_), .Q(reg_pc_21_) );
DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf112), .D(_84__22_), .Q(reg_pc_22_) );
DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf111), .D(_84__23_), .Q(reg_pc_23_) );
DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf110), .D(_84__24_), .Q(reg_pc_24_) );
DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf109), .D(_84__25_), .Q(reg_pc_25_) );
DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf108), .D(_84__26_), .Q(reg_pc_26_) );
DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf107), .D(_84__27_), .Q(reg_pc_27_) );
DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf106), .D(_84__28_), .Q(reg_pc_28_) );
DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf105), .D(_84__29_), .Q(reg_pc_29_) );
DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf104), .D(_84__30_), .Q(reg_pc_30_) );
DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf103), .D(_84__31_), .Q(reg_pc_31_) );
DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf102), .D(_80__0_), .Q(reg_next_pc_0_) );
DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf101), .D(_80__1_), .Q(reg_next_pc_1_) );
DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf100), .D(_80__2_), .Q(reg_next_pc_2_) );
DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf99), .D(_80__3_), .Q(reg_next_pc_3_) );
DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf98), .D(_80__4_), .Q(reg_next_pc_4_) );
DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf97), .D(_80__5_), .Q(reg_next_pc_5_) );
DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf96), .D(_80__6_), .Q(reg_next_pc_6_) );
DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf95), .D(_80__7_), .Q(reg_next_pc_7_) );
DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf94), .D(_80__8_), .Q(reg_next_pc_8_) );
DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf93), .D(_80__9_), .Q(reg_next_pc_9_) );
DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf92), .D(_80__10_), .Q(reg_next_pc_10_) );
DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf91), .D(_80__11_), .Q(reg_next_pc_11_) );
DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf90), .D(_80__12_), .Q(reg_next_pc_12_) );
DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf89), .D(_80__13_), .Q(reg_next_pc_13_) );
DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf88), .D(_80__14_), .Q(reg_next_pc_14_) );
DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf87), .D(_80__15_), .Q(reg_next_pc_15_) );
DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf86), .D(_80__16_), .Q(reg_next_pc_16_) );
DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf85), .D(_80__17_), .Q(reg_next_pc_17_) );
DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf84), .D(_80__18_), .Q(reg_next_pc_18_) );
DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf83), .D(_80__19_), .Q(reg_next_pc_19_) );
DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf82), .D(_80__20_), .Q(reg_next_pc_20_) );
DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf81), .D(_80__21_), .Q(reg_next_pc_21_) );
DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf80), .D(_80__22_), .Q(reg_next_pc_22_) );
DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf79), .D(_80__23_), .Q(reg_next_pc_23_) );
DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf78), .D(_80__24_), .Q(reg_next_pc_24_) );
DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf77), .D(_80__25_), .Q(reg_next_pc_25_) );
DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf76), .D(_80__26_), .Q(reg_next_pc_26_) );
DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf75), .D(_80__27_), .Q(reg_next_pc_27_) );
DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf74), .D(_80__28_), .Q(reg_next_pc_28_) );
DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf73), .D(_80__29_), .Q(reg_next_pc_29_) );
DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf72), .D(_80__30_), .Q(reg_next_pc_30_) );
DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf71), .D(_80__31_), .Q(reg_next_pc_31_) );
DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf70), .D(_81__0_), .Q(_10734__0_) );
DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf69), .D(_81__1_), .Q(_10734__1_) );
DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf68), .D(_81__2_), .Q(_10734__2_) );
DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf67), .D(_81__3_), .Q(_10734__3_) );
DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf66), .D(_81__4_), .Q(_10734__4_) );
DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf65), .D(_81__5_), .Q(_10734__5_) );
DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf64), .D(_81__6_), .Q(_10734__6_) );
DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf63), .D(_81__7_), .Q(_10734__7_) );
DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf62), .D(_81__8_), .Q(_10734__8_) );
DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf61), .D(_81__9_), .Q(_10734__9_) );
DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf60), .D(_81__10_), .Q(_10734__10_) );
DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf59), .D(_81__11_), .Q(_10734__11_) );
DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf58), .D(_81__12_), .Q(_10734__12_) );
DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf57), .D(_81__13_), .Q(_10734__13_) );
DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf56), .D(_81__14_), .Q(_10734__14_) );
DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf55), .D(_81__15_), .Q(_10734__15_) );
DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf54), .D(_81__16_), .Q(_10734__16_) );
DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf53), .D(_81__17_), .Q(_10734__17_) );
DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf52), .D(_81__18_), .Q(_10734__18_) );
DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf51), .D(_81__19_), .Q(_10734__19_) );
DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf50), .D(_81__20_), .Q(_10734__20_) );
DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf49), .D(_81__21_), .Q(_10734__21_) );
DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf48), .D(_81__22_), .Q(_10734__22_) );
DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf47), .D(_81__23_), .Q(_10734__23_) );
DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf46), .D(_81__24_), .Q(_10734__24_) );
DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf45), .D(_81__25_), .Q(_10734__25_) );
DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf44), .D(_81__26_), .Q(_10734__26_) );
DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf43), .D(_81__27_), .Q(_10734__27_) );
DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf42), .D(_81__28_), .Q(_10734__28_) );
DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf41), .D(_81__29_), .Q(_10734__29_) );
DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf40), .D(_81__30_), .Q(_10734__30_) );
DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf39), .D(_81__31_), .Q(_10734__31_) );
DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf38), .D(_82__0_), .Q(_10728__0_) );
DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf37), .D(_82__1_), .Q(_10728__1_) );
DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf36), .D(_82__2_), .Q(_10728__2_) );
DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf35), .D(_82__3_), .Q(_10728__3_) );
DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf34), .D(_82__4_), .Q(_10728__4_) );
DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf33), .D(_82__5_), .Q(_10728__5_) );
DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf32), .D(_82__6_), .Q(_10728__6_) );
DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf31), .D(_82__7_), .Q(_10728__7_) );
DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf30), .D(_82__8_), .Q(_10735__8_) );
DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf29), .D(_82__9_), .Q(_10735__9_) );
DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf28), .D(_82__10_), .Q(_10735__10_) );
DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf27), .D(_82__11_), .Q(_10735__11_) );
DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf26), .D(_82__12_), .Q(_10735__12_) );
DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf25), .D(_82__13_), .Q(_10735__13_) );
DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf24), .D(_82__14_), .Q(_10735__14_) );
DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf23), .D(_82__15_), .Q(_10735__15_) );
DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf22), .D(_82__16_), .Q(_10735__16_) );
DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf21), .D(_82__17_), .Q(_10735__17_) );
DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf20), .D(_82__18_), .Q(_10735__18_) );
DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf19), .D(_82__19_), .Q(_10735__19_) );
DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf18), .D(_82__20_), .Q(_10735__20_) );
DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf17), .D(_82__21_), .Q(_10735__21_) );
DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf16), .D(_82__22_), .Q(_10735__22_) );
DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf15), .D(_82__23_), .Q(_10735__23_) );
DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf14), .D(_82__24_), .Q(_10735__24_) );
DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf13), .D(_82__25_), .Q(_10735__25_) );
DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf12), .D(_82__26_), .Q(_10735__26_) );
DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf11), .D(_82__27_), .Q(_10735__27_) );
DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf10), .D(_82__28_), .Q(_10735__28_) );
DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf9), .D(_82__29_), .Q(_10735__29_) );
DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf8), .D(_82__30_), .Q(_10735__30_) );
DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf7), .D(_82__31_), .Q(_10735__31_) );
DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf6), .D(_83__0_), .Q(reg_out_0_) );
DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf5), .D(_83__1_), .Q(reg_out_1_) );
DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf4), .D(_83__2_), .Q(reg_out_2_) );
DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf3), .D(_83__3_), .Q(reg_out_3_) );
DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf2), .D(_83__4_), .Q(reg_out_4_) );
DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf1), .D(_83__5_), .Q(reg_out_5_) );
DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf0), .D(_83__6_), .Q(reg_out_6_) );
DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf136), .D(_83__7_), .Q(reg_out_7_) );
DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf135), .D(_83__8_), .Q(reg_out_8_) );
DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf134), .D(_83__9_), .Q(reg_out_9_) );
DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf133), .D(_83__10_), .Q(reg_out_10_) );
DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf132), .D(_83__11_), .Q(reg_out_11_) );
DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf131), .D(_83__12_), .Q(reg_out_12_) );
DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf130), .D(_83__13_), .Q(reg_out_13_) );
DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf129), .D(_83__14_), .Q(reg_out_14_) );
DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf128), .D(_83__15_), .Q(reg_out_15_) );
DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf127), .D(_83__16_), .Q(reg_out_16_) );
DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf126), .D(_83__17_), .Q(reg_out_17_) );
DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf125), .D(_83__18_), .Q(reg_out_18_) );
DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf124), .D(_83__19_), .Q(reg_out_19_) );
DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf123), .D(_83__20_), .Q(reg_out_20_) );
DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf122), .D(_83__21_), .Q(reg_out_21_) );
DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf121), .D(_83__22_), .Q(reg_out_22_) );
DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf120), .D(_83__23_), .Q(reg_out_23_) );
DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf119), .D(_83__24_), .Q(reg_out_24_) );
DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf118), .D(_83__25_), .Q(reg_out_25_) );
DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf117), .D(_83__26_), .Q(reg_out_26_) );
DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf116), .D(_83__27_), .Q(reg_out_27_) );
DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf115), .D(_83__28_), .Q(reg_out_28_) );
DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf114), .D(_83__29_), .Q(reg_out_29_) );
DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf113), .D(_83__30_), .Q(reg_out_30_) );
DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf112), .D(_83__31_), .Q(reg_out_31_) );
DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf111), .D(_85__0_), .Q(reg_sh_0_) );
DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf110), .D(_85__1_), .Q(reg_sh_1_) );
DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf109), .D(_85__2_), .Q(reg_sh_2_) );
DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf108), .D(_85__3_), .Q(reg_sh_3_) );
DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf107), .D(_85__4_), .Q(reg_sh_4_) );
DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf106), .D(_71_), .Q(mem_do_prefetch) );
DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf105), .D(_73_), .Q(mem_do_rinst) );
DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf104), .D(_72_), .Q(mem_do_rdata) );
DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf103), .D(_74_), .Q(mem_do_wdata) );
DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf102), .D(_8_), .Q(decoder_trigger) );
DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf101), .D(_7_), .Q(decoder_pseudo_trigger) );
DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf100), .D(_69_), .Q(latched_store) );
DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf99), .D(_68_), .Q(latched_stalu) );
DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf98), .D(_63_), .Q(latched_branch) );
DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf97), .D(_64_), .Q(latched_compr) );
DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf96), .D(_66_), .Q(latched_is_lu) );
DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf95), .D(_65_), .Q(latched_is_lh) );
DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf94), .D(_67__0_), .Q(latched_rd_0_) );
DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf93), .D(_67__1_), .Q(latched_rd_1_) );
DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf92), .D(_67__2_), .Q(latched_rd_2_) );
DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf91), .D(_67__3_), .Q(latched_rd_3_) );
DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf90), .D(_67__4_), .Q(latched_rd_4_) );
DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf89), .D(alu_out_0_), .Q(alu_out_q_0_) );
DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf88), .D(alu_out_1_), .Q(alu_out_q_1_) );
DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf87), .D(alu_out_2_), .Q(alu_out_q_2_) );
DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf86), .D(alu_out_3_), .Q(alu_out_q_3_) );
DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf85), .D(alu_out_4_), .Q(alu_out_q_4_) );
DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf84), .D(alu_out_5_), .Q(alu_out_q_5_) );
DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf83), .D(alu_out_6_), .Q(alu_out_q_6_) );
DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf82), .D(alu_out_7_), .Q(alu_out_q_7_) );
DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf81), .D(alu_out_8_), .Q(alu_out_q_8_) );
DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf80), .D(alu_out_9_), .Q(alu_out_q_9_) );
DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf79), .D(alu_out_10_), .Q(alu_out_q_10_) );
DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf78), .D(alu_out_11_), .Q(alu_out_q_11_) );
DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf77), .D(alu_out_12_), .Q(alu_out_q_12_) );
DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf76), .D(alu_out_13_), .Q(alu_out_q_13_) );
DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf75), .D(alu_out_14_), .Q(alu_out_q_14_) );
DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf74), .D(alu_out_15_), .Q(alu_out_q_15_) );
DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf73), .D(alu_out_16_), .Q(alu_out_q_16_) );
DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf72), .D(alu_out_17_), .Q(alu_out_q_17_) );
DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf71), .D(alu_out_18_), .Q(alu_out_q_18_) );
DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf70), .D(alu_out_19_), .Q(alu_out_q_19_) );
DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf69), .D(alu_out_20_), .Q(alu_out_q_20_) );
DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf68), .D(alu_out_21_), .Q(alu_out_q_21_) );
DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf67), .D(alu_out_22_), .Q(alu_out_q_22_) );
DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf66), .D(alu_out_23_), .Q(alu_out_q_23_) );
DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf65), .D(alu_out_24_), .Q(alu_out_q_24_) );
DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf64), .D(alu_out_25_), .Q(alu_out_q_25_) );
DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf63), .D(alu_out_26_), .Q(alu_out_q_26_) );
DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf62), .D(alu_out_27_), .Q(alu_out_q_27_) );
DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf61), .D(alu_out_28_), .Q(alu_out_q_28_) );
DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf60), .D(alu_out_29_), .Q(alu_out_q_29_) );
DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf59), .D(alu_out_30_), .Q(alu_out_q_30_) );
DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf58), .D(alu_out_31_), .Q(alu_out_q_31_) );
DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf57), .D(_26_), .Q(instr_lui) );
DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf56), .D(_13_), .Q(instr_auipc) );
DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf55), .D(_20_), .Q(instr_jal) );
DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf54), .D(_21_), .Q(instr_jalr) );
DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf53), .D(_14_), .Q(instr_beq) );
DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf52), .D(_19_), .Q(instr_bne) );
DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf51), .D(_17_), .Q(instr_blt) );
DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf50), .D(_15_), .Q(instr_bge) );
DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf49), .D(_18_), .Q(instr_bltu) );
DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf48), .D(_16_), .Q(instr_bgeu) );
DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf47), .D(_22_), .Q(instr_lb) );
DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf46), .D(_24_), .Q(instr_lh) );
DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf45), .D(_27_), .Q(instr_lw) );
DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf44), .D(_23_), .Q(instr_lbu) );
DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf43), .D(_25_), .Q(instr_lhu) );
DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf42), .D(_34_), .Q(instr_sb) );
DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf41), .D(_35_), .Q(instr_sh) );
DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf40), .D(_47_), .Q(instr_sw) );
DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf39), .D(_10_), .Q(instr_addi) );
DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf38), .D(_39_), .Q(instr_slti) );
DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf37), .D(_40_), .Q(instr_sltiu) );
DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf36), .D(_49_), .Q(instr_xori) );
DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf35), .D(_29_), .Q(instr_ori) );
DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf34), .D(_12_), .Q(instr_andi) );
DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf33), .D(_37_), .Q(instr_slli) );
DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf32), .D(_45_), .Q(instr_srli) );
DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf31), .D(_43_), .Q(instr_srai) );
DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf30), .D(_9_), .Q(instr_add) );
DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf29), .D(_46_), .Q(instr_sub) );
DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf28), .D(_36_), .Q(instr_sll) );
DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_bF_buf27), .D(_38_), .Q(instr_slt) );
DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_bF_buf26), .D(_41_), .Q(instr_sltu) );
DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_bF_buf25), .D(_48_), .Q(instr_xor) );
DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_bF_buf24), .D(_44_), .Q(instr_srl) );
DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_bF_buf23), .D(_42_), .Q(instr_sra) );
DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_bF_buf22), .D(_28_), .Q(instr_or) );
DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_bF_buf21), .D(_11_), .Q(instr_and) );
DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_bF_buf20), .D(_30_), .Q(instr_rdcycle) );
DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_bF_buf19), .D(_31_), .Q(instr_rdcycleh) );
DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_bF_buf18), .D(_32_), .Q(instr_rdinstr) );
DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_bF_buf17), .D(_33_), .Q(instr_rdinstrh) );
DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_bF_buf16), .D(_4__0_), .Q(decoded_rd_0_) );
DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_bF_buf15), .D(_4__1_), .Q(decoded_rd_1_) );
DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_bF_buf14), .D(_4__2_), .Q(decoded_rd_2_) );
DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_bF_buf13), .D(_4__3_), .Q(decoded_rd_3_) );
DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_bF_buf12), .D(_4__4_), .Q(decoded_rd_4_) );
DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_bF_buf11), .D(_2__0_), .Q(decoded_imm_0_) );
DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_bF_buf10), .D(_2__1_), .Q(decoded_imm_1_) );
DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_bF_buf9), .D(_2__2_), .Q(decoded_imm_2_) );
DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_bF_buf8), .D(_2__3_), .Q(decoded_imm_3_) );
DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_bF_buf7), .D(_2__4_), .Q(decoded_imm_4_) );
DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_bF_buf6), .D(_2__5_), .Q(decoded_imm_5_) );
DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_bF_buf5), .D(_2__6_), .Q(decoded_imm_6_) );
DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_bF_buf4), .D(_2__7_), .Q(decoded_imm_7_) );
DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_bF_buf3), .D(_2__8_), .Q(decoded_imm_8_) );
DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_bF_buf2), .D(_2__9_), .Q(decoded_imm_9_) );
DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_bF_buf1), .D(_2__10_), .Q(decoded_imm_10_) );
DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_bF_buf0), .D(_2__11_), .Q(decoded_imm_11_) );
DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_bF_buf136), .D(_2__12_), .Q(decoded_imm_12_) );
DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_bF_buf135), .D(_2__13_), .Q(decoded_imm_13_) );
DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_bF_buf134), .D(_2__14_), .Q(decoded_imm_14_) );
DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_bF_buf133), .D(_2__15_), .Q(decoded_imm_15_) );
DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_bF_buf132), .D(_2__16_), .Q(decoded_imm_16_) );
DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_bF_buf131), .D(_2__17_), .Q(decoded_imm_17_) );
DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_bF_buf130), .D(_2__18_), .Q(decoded_imm_18_) );
DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_bF_buf129), .D(_2__19_), .Q(decoded_imm_19_) );
DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_bF_buf128), .D(_2__20_), .Q(decoded_imm_20_) );
DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_bF_buf127), .D(_2__21_), .Q(decoded_imm_21_) );
DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_bF_buf126), .D(_2__22_), .Q(decoded_imm_22_) );
DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_bF_buf125), .D(_2__23_), .Q(decoded_imm_23_) );
DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_bF_buf124), .D(_2__24_), .Q(decoded_imm_24_) );
DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_bF_buf123), .D(_2__25_), .Q(decoded_imm_25_) );
DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_bF_buf122), .D(_2__26_), .Q(decoded_imm_26_) );
DFFPOSX1 DFFPOSX1_838 ( .CLK(clk_bF_buf121), .D(_2__27_), .Q(decoded_imm_27_) );
DFFPOSX1 DFFPOSX1_839 ( .CLK(clk_bF_buf120), .D(_2__28_), .Q(decoded_imm_28_) );
DFFPOSX1 DFFPOSX1_840 ( .CLK(clk_bF_buf119), .D(_2__29_), .Q(decoded_imm_29_) );
DFFPOSX1 DFFPOSX1_841 ( .CLK(clk_bF_buf118), .D(_2__30_), .Q(decoded_imm_30_) );
DFFPOSX1 DFFPOSX1_842 ( .CLK(clk_bF_buf117), .D(_2__31_), .Q(decoded_imm_31_) );
DFFPOSX1 DFFPOSX1_843 ( .CLK(clk_bF_buf116), .D(_3__0_), .Q(decoded_imm_uj_0_) );
DFFPOSX1 DFFPOSX1_844 ( .CLK(clk_bF_buf115), .D(_3__1_), .Q(decoded_imm_uj_1_) );
DFFPOSX1 DFFPOSX1_845 ( .CLK(clk_bF_buf114), .D(_3__2_), .Q(decoded_imm_uj_2_) );
DFFPOSX1 DFFPOSX1_846 ( .CLK(clk_bF_buf113), .D(_3__3_), .Q(decoded_imm_uj_3_) );
DFFPOSX1 DFFPOSX1_847 ( .CLK(clk_bF_buf112), .D(_3__4_), .Q(decoded_imm_uj_4_) );
DFFPOSX1 DFFPOSX1_848 ( .CLK(clk_bF_buf111), .D(_3__5_), .Q(decoded_imm_uj_5_) );
DFFPOSX1 DFFPOSX1_849 ( .CLK(clk_bF_buf110), .D(_3__6_), .Q(decoded_imm_uj_6_) );
DFFPOSX1 DFFPOSX1_850 ( .CLK(clk_bF_buf109), .D(_3__7_), .Q(decoded_imm_uj_7_) );
DFFPOSX1 DFFPOSX1_851 ( .CLK(clk_bF_buf108), .D(_3__8_), .Q(decoded_imm_uj_8_) );
DFFPOSX1 DFFPOSX1_852 ( .CLK(clk_bF_buf107), .D(_3__9_), .Q(decoded_imm_uj_9_) );
DFFPOSX1 DFFPOSX1_853 ( .CLK(clk_bF_buf106), .D(_3__10_), .Q(decoded_imm_uj_10_) );
DFFPOSX1 DFFPOSX1_854 ( .CLK(clk_bF_buf105), .D(_3__11_), .Q(decoded_imm_uj_11_) );
DFFPOSX1 DFFPOSX1_855 ( .CLK(clk_bF_buf104), .D(_3__12_), .Q(decoded_imm_uj_12_) );
DFFPOSX1 DFFPOSX1_856 ( .CLK(clk_bF_buf103), .D(_3__13_), .Q(decoded_imm_uj_13_) );
DFFPOSX1 DFFPOSX1_857 ( .CLK(clk_bF_buf102), .D(_3__14_), .Q(decoded_imm_uj_14_) );
DFFPOSX1 DFFPOSX1_858 ( .CLK(clk_bF_buf101), .D(_3__15_), .Q(decoded_imm_uj_15_) );
DFFPOSX1 DFFPOSX1_859 ( .CLK(clk_bF_buf100), .D(_3__16_), .Q(decoded_imm_uj_16_) );
DFFPOSX1 DFFPOSX1_860 ( .CLK(clk_bF_buf99), .D(_3__17_), .Q(decoded_imm_uj_17_) );
DFFPOSX1 DFFPOSX1_861 ( .CLK(clk_bF_buf98), .D(_3__18_), .Q(decoded_imm_uj_18_) );
DFFPOSX1 DFFPOSX1_862 ( .CLK(clk_bF_buf97), .D(_3__19_), .Q(decoded_imm_uj_19_) );
DFFPOSX1 DFFPOSX1_863 ( .CLK(clk_bF_buf96), .D(_3__20_), .Q(decoded_imm_uj_20_) );
DFFPOSX1 DFFPOSX1_864 ( .CLK(clk_bF_buf95), .D(_3__21_), .Q(decoded_imm_uj_21_) );
DFFPOSX1 DFFPOSX1_865 ( .CLK(clk_bF_buf94), .D(_3__22_), .Q(decoded_imm_uj_22_) );
DFFPOSX1 DFFPOSX1_866 ( .CLK(clk_bF_buf93), .D(_3__23_), .Q(decoded_imm_uj_23_) );
DFFPOSX1 DFFPOSX1_867 ( .CLK(clk_bF_buf92), .D(_3__24_), .Q(decoded_imm_uj_24_) );
DFFPOSX1 DFFPOSX1_868 ( .CLK(clk_bF_buf91), .D(_3__25_), .Q(decoded_imm_uj_25_) );
DFFPOSX1 DFFPOSX1_869 ( .CLK(clk_bF_buf90), .D(_3__26_), .Q(decoded_imm_uj_26_) );
DFFPOSX1 DFFPOSX1_870 ( .CLK(clk_bF_buf89), .D(_3__27_), .Q(decoded_imm_uj_27_) );
DFFPOSX1 DFFPOSX1_871 ( .CLK(clk_bF_buf88), .D(_3__28_), .Q(decoded_imm_uj_28_) );
DFFPOSX1 DFFPOSX1_872 ( .CLK(clk_bF_buf87), .D(_3__29_), .Q(decoded_imm_uj_29_) );
DFFPOSX1 DFFPOSX1_873 ( .CLK(clk_bF_buf86), .D(_3__30_), .Q(decoded_imm_uj_30_) );
DFFPOSX1 DFFPOSX1_874 ( .CLK(clk_bF_buf85), .D(_3__31_), .Q(decoded_imm_uj_31_) );
DFFPOSX1 DFFPOSX1_875 ( .CLK(clk_bF_buf84), .D(_57_), .Q(is_lui_auipc_jal) );
DFFPOSX1 DFFPOSX1_876 ( .CLK(clk_bF_buf83), .D(_55_), .Q(is_lb_lh_lw_lbu_lhu) );
DFFPOSX1 DFFPOSX1_877 ( .CLK(clk_bF_buf82), .D(_61_), .Q(is_slli_srli_srai) );
DFFPOSX1 DFFPOSX1_878 ( .CLK(clk_bF_buf81), .D(_54_), .Q(is_jalr_addi_slti_sltiu_xori_ori_andi) );
DFFPOSX1 DFFPOSX1_879 ( .CLK(clk_bF_buf80), .D(_59_), .Q(is_sb_sh_sw) );
DFFPOSX1 DFFPOSX1_880 ( .CLK(clk_bF_buf79), .D(_60_), .Q(is_sll_srl_sra) );
DFFPOSX1 DFFPOSX1_881 ( .CLK(clk_bF_buf78), .D(_58_), .Q(is_lui_auipc_jal_jalr_addi_add_sub) );
DFFPOSX1 DFFPOSX1_882 ( .CLK(clk_bF_buf77), .D(_62_), .Q(is_slti_blt_slt) );
DFFPOSX1 DFFPOSX1_883 ( .CLK(clk_bF_buf76), .D(_52_), .Q(is_beq_bne_blt_bge_bltu_bgeu) );
DFFPOSX1 DFFPOSX1_884 ( .CLK(clk_bF_buf75), .D(_56_), .Q(is_lbu_lhu_lw) );
DFFPOSX1 DFFPOSX1_885 ( .CLK(clk_bF_buf74), .D(_50_), .Q(is_alu_reg_imm) );
DFFPOSX1 DFFPOSX1_886 ( .CLK(clk_bF_buf73), .D(_51_), .Q(is_alu_reg_reg) );
DFFPOSX1 DFFPOSX1_887 ( .CLK(clk_bF_buf72), .D(_53_), .Q(is_compare) );
DFFPOSX1 DFFPOSX1_888 ( .CLK(clk_bF_buf71), .D(_77_), .Q(_10731_) );
DFFPOSX1 DFFPOSX1_889 ( .CLK(clk_bF_buf70), .D(_75_), .Q(_10725_) );
DFFPOSX1 DFFPOSX1_890 ( .CLK(clk_bF_buf69), .D(_70__0_), .Q(_10724__0_) );
DFFPOSX1 DFFPOSX1_891 ( .CLK(clk_bF_buf68), .D(_70__1_), .Q(_10724__1_) );
DFFPOSX1 DFFPOSX1_892 ( .CLK(clk_bF_buf67), .D(_70__2_), .Q(_10724__2_) );
DFFPOSX1 DFFPOSX1_893 ( .CLK(clk_bF_buf66), .D(_70__3_), .Q(_10724__3_) );
DFFPOSX1 DFFPOSX1_894 ( .CLK(clk_bF_buf65), .D(_70__4_), .Q(_10724__4_) );
DFFPOSX1 DFFPOSX1_895 ( .CLK(clk_bF_buf64), .D(_70__5_), .Q(_10724__5_) );
DFFPOSX1 DFFPOSX1_896 ( .CLK(clk_bF_buf63), .D(_70__6_), .Q(_10724__6_) );
DFFPOSX1 DFFPOSX1_897 ( .CLK(clk_bF_buf62), .D(_70__7_), .Q(_10724__7_) );
DFFPOSX1 DFFPOSX1_898 ( .CLK(clk_bF_buf61), .D(_70__8_), .Q(_10724__8_) );
DFFPOSX1 DFFPOSX1_899 ( .CLK(clk_bF_buf60), .D(_70__9_), .Q(_10724__9_) );
DFFPOSX1 DFFPOSX1_900 ( .CLK(clk_bF_buf59), .D(_70__10_), .Q(_10724__10_) );
DFFPOSX1 DFFPOSX1_901 ( .CLK(clk_bF_buf58), .D(_70__11_), .Q(_10724__11_) );
DFFPOSX1 DFFPOSX1_902 ( .CLK(clk_bF_buf57), .D(_70__12_), .Q(_10724__12_) );
DFFPOSX1 DFFPOSX1_903 ( .CLK(clk_bF_buf56), .D(_70__13_), .Q(_10724__13_) );
DFFPOSX1 DFFPOSX1_904 ( .CLK(clk_bF_buf55), .D(_70__14_), .Q(_10724__14_) );
DFFPOSX1 DFFPOSX1_905 ( .CLK(clk_bF_buf54), .D(_70__15_), .Q(_10724__15_) );
DFFPOSX1 DFFPOSX1_906 ( .CLK(clk_bF_buf53), .D(_70__16_), .Q(_10724__16_) );
DFFPOSX1 DFFPOSX1_907 ( .CLK(clk_bF_buf52), .D(_70__17_), .Q(_10724__17_) );
DFFPOSX1 DFFPOSX1_908 ( .CLK(clk_bF_buf51), .D(_70__18_), .Q(_10724__18_) );
DFFPOSX1 DFFPOSX1_909 ( .CLK(clk_bF_buf50), .D(_70__19_), .Q(_10724__19_) );
DFFPOSX1 DFFPOSX1_910 ( .CLK(clk_bF_buf49), .D(_70__20_), .Q(_10724__20_) );
DFFPOSX1 DFFPOSX1_911 ( .CLK(clk_bF_buf48), .D(_70__21_), .Q(_10724__21_) );
DFFPOSX1 DFFPOSX1_912 ( .CLK(clk_bF_buf47), .D(_70__22_), .Q(_10724__22_) );
DFFPOSX1 DFFPOSX1_913 ( .CLK(clk_bF_buf46), .D(_70__23_), .Q(_10724__23_) );
DFFPOSX1 DFFPOSX1_914 ( .CLK(clk_bF_buf45), .D(_70__24_), .Q(_10724__24_) );
DFFPOSX1 DFFPOSX1_915 ( .CLK(clk_bF_buf44), .D(_70__25_), .Q(_10724__25_) );
DFFPOSX1 DFFPOSX1_916 ( .CLK(clk_bF_buf43), .D(_70__26_), .Q(_10724__26_) );
DFFPOSX1 DFFPOSX1_917 ( .CLK(clk_bF_buf42), .D(_70__27_), .Q(_10724__27_) );
DFFPOSX1 DFFPOSX1_918 ( .CLK(clk_bF_buf41), .D(_70__28_), .Q(_10724__28_) );
DFFPOSX1 DFFPOSX1_919 ( .CLK(clk_bF_buf40), .D(_70__29_), .Q(_10724__29_) );
DFFPOSX1 DFFPOSX1_920 ( .CLK(clk_bF_buf39), .D(_70__30_), .Q(_10724__30_) );
DFFPOSX1 DFFPOSX1_921 ( .CLK(clk_bF_buf38), .D(_70__31_), .Q(_10724__31_) );
DFFPOSX1 DFFPOSX1_922 ( .CLK(clk_bF_buf37), .D(_78__0_), .Q(_10732__0_) );
DFFPOSX1 DFFPOSX1_923 ( .CLK(clk_bF_buf36), .D(_78__1_), .Q(_10732__1_) );
DFFPOSX1 DFFPOSX1_924 ( .CLK(clk_bF_buf35), .D(_78__2_), .Q(_10732__2_) );
DFFPOSX1 DFFPOSX1_925 ( .CLK(clk_bF_buf34), .D(_78__3_), .Q(_10732__3_) );
DFFPOSX1 DFFPOSX1_926 ( .CLK(clk_bF_buf33), .D(_78__4_), .Q(_10732__4_) );
DFFPOSX1 DFFPOSX1_927 ( .CLK(clk_bF_buf32), .D(_78__5_), .Q(_10732__5_) );
DFFPOSX1 DFFPOSX1_928 ( .CLK(clk_bF_buf31), .D(_78__6_), .Q(_10732__6_) );
DFFPOSX1 DFFPOSX1_929 ( .CLK(clk_bF_buf30), .D(_78__7_), .Q(_10732__7_) );
DFFPOSX1 DFFPOSX1_930 ( .CLK(clk_bF_buf29), .D(_78__8_), .Q(_10732__8_) );
DFFPOSX1 DFFPOSX1_931 ( .CLK(clk_bF_buf28), .D(_78__9_), .Q(_10732__9_) );
DFFPOSX1 DFFPOSX1_932 ( .CLK(clk_bF_buf27), .D(_78__10_), .Q(_10732__10_) );
DFFPOSX1 DFFPOSX1_933 ( .CLK(clk_bF_buf26), .D(_78__11_), .Q(_10732__11_) );
DFFPOSX1 DFFPOSX1_934 ( .CLK(clk_bF_buf25), .D(_78__12_), .Q(_10732__12_) );
DFFPOSX1 DFFPOSX1_935 ( .CLK(clk_bF_buf24), .D(_78__13_), .Q(_10732__13_) );
DFFPOSX1 DFFPOSX1_936 ( .CLK(clk_bF_buf23), .D(_78__14_), .Q(_10732__14_) );
DFFPOSX1 DFFPOSX1_937 ( .CLK(clk_bF_buf22), .D(_78__15_), .Q(_10732__15_) );
DFFPOSX1 DFFPOSX1_938 ( .CLK(clk_bF_buf21), .D(_78__16_), .Q(_10732__16_) );
DFFPOSX1 DFFPOSX1_939 ( .CLK(clk_bF_buf20), .D(_78__17_), .Q(_10732__17_) );
DFFPOSX1 DFFPOSX1_940 ( .CLK(clk_bF_buf19), .D(_78__18_), .Q(_10732__18_) );
DFFPOSX1 DFFPOSX1_941 ( .CLK(clk_bF_buf18), .D(_78__19_), .Q(_10732__19_) );
DFFPOSX1 DFFPOSX1_942 ( .CLK(clk_bF_buf17), .D(_78__20_), .Q(_10732__20_) );
DFFPOSX1 DFFPOSX1_943 ( .CLK(clk_bF_buf16), .D(_78__21_), .Q(_10732__21_) );
DFFPOSX1 DFFPOSX1_944 ( .CLK(clk_bF_buf15), .D(_78__22_), .Q(_10732__22_) );
DFFPOSX1 DFFPOSX1_945 ( .CLK(clk_bF_buf14), .D(_78__23_), .Q(_10732__23_) );
DFFPOSX1 DFFPOSX1_946 ( .CLK(clk_bF_buf13), .D(_78__24_), .Q(_10732__24_) );
DFFPOSX1 DFFPOSX1_947 ( .CLK(clk_bF_buf12), .D(_78__25_), .Q(_10732__25_) );
DFFPOSX1 DFFPOSX1_948 ( .CLK(clk_bF_buf11), .D(_78__26_), .Q(_10732__26_) );
DFFPOSX1 DFFPOSX1_949 ( .CLK(clk_bF_buf10), .D(_78__27_), .Q(_10732__27_) );
DFFPOSX1 DFFPOSX1_950 ( .CLK(clk_bF_buf9), .D(_78__28_), .Q(_10732__28_) );
DFFPOSX1 DFFPOSX1_951 ( .CLK(clk_bF_buf8), .D(_78__29_), .Q(_10732__29_) );
DFFPOSX1 DFFPOSX1_952 ( .CLK(clk_bF_buf7), .D(_78__30_), .Q(_10732__30_) );
DFFPOSX1 DFFPOSX1_953 ( .CLK(clk_bF_buf6), .D(_78__31_), .Q(_10732__31_) );
DFFPOSX1 DFFPOSX1_954 ( .CLK(clk_bF_buf5), .D(_79__0_), .Q(_10733__0_) );
DFFPOSX1 DFFPOSX1_955 ( .CLK(clk_bF_buf4), .D(_79__1_), .Q(_10733__1_) );
DFFPOSX1 DFFPOSX1_956 ( .CLK(clk_bF_buf3), .D(_79__2_), .Q(_10733__2_) );
DFFPOSX1 DFFPOSX1_957 ( .CLK(clk_bF_buf2), .D(_79__3_), .Q(_10733__3_) );
DFFPOSX1 DFFPOSX1_958 ( .CLK(clk_bF_buf1), .D(_76__0_), .Q(mem_state_0_) );
DFFPOSX1 DFFPOSX1_959 ( .CLK(clk_bF_buf0), .D(_76__1_), .Q(mem_state_1_) );
DFFPOSX1 DFFPOSX1_960 ( .CLK(clk_bF_buf136), .D(mem_rdata_latched_0_), .Q(mem_rdata_q_0_) );
DFFPOSX1 DFFPOSX1_961 ( .CLK(clk_bF_buf135), .D(mem_rdata_latched_1_), .Q(mem_rdata_q_1_) );
DFFPOSX1 DFFPOSX1_962 ( .CLK(clk_bF_buf134), .D(mem_rdata_latched_2_), .Q(mem_rdata_q_2_) );
DFFPOSX1 DFFPOSX1_963 ( .CLK(clk_bF_buf133), .D(mem_rdata_latched_3_), .Q(mem_rdata_q_3_) );
DFFPOSX1 DFFPOSX1_964 ( .CLK(clk_bF_buf132), .D(mem_rdata_latched_4_), .Q(mem_rdata_q_4_) );
DFFPOSX1 DFFPOSX1_965 ( .CLK(clk_bF_buf131), .D(mem_rdata_latched_5_), .Q(mem_rdata_q_5_) );
DFFPOSX1 DFFPOSX1_966 ( .CLK(clk_bF_buf130), .D(mem_rdata_latched_6_), .Q(mem_rdata_q_6_) );
DFFPOSX1 DFFPOSX1_967 ( .CLK(clk_bF_buf129), .D(mem_rdata_latched_7_), .Q(mem_rdata_q_7_) );
DFFPOSX1 DFFPOSX1_968 ( .CLK(clk_bF_buf128), .D(mem_rdata_latched_8_), .Q(mem_rdata_q_8_) );
DFFPOSX1 DFFPOSX1_969 ( .CLK(clk_bF_buf127), .D(mem_rdata_latched_9_), .Q(mem_rdata_q_9_) );
DFFPOSX1 DFFPOSX1_970 ( .CLK(clk_bF_buf126), .D(mem_rdata_latched_10_), .Q(mem_rdata_q_10_) );
DFFPOSX1 DFFPOSX1_971 ( .CLK(clk_bF_buf125), .D(mem_rdata_latched_11_), .Q(mem_rdata_q_11_) );
DFFPOSX1 DFFPOSX1_972 ( .CLK(clk_bF_buf124), .D(mem_rdata_latched_12_), .Q(mem_rdata_q_12_) );
DFFPOSX1 DFFPOSX1_973 ( .CLK(clk_bF_buf123), .D(mem_rdata_latched_13_), .Q(mem_rdata_q_13_) );
DFFPOSX1 DFFPOSX1_974 ( .CLK(clk_bF_buf122), .D(mem_rdata_latched_14_), .Q(mem_rdata_q_14_) );
DFFPOSX1 DFFPOSX1_975 ( .CLK(clk_bF_buf121), .D(mem_rdata_latched_15_), .Q(mem_rdata_q_15_) );
DFFPOSX1 DFFPOSX1_976 ( .CLK(clk_bF_buf120), .D(mem_rdata_latched_16_), .Q(mem_rdata_q_16_) );
DFFPOSX1 DFFPOSX1_977 ( .CLK(clk_bF_buf119), .D(mem_rdata_latched_17_), .Q(mem_rdata_q_17_) );
DFFPOSX1 DFFPOSX1_978 ( .CLK(clk_bF_buf118), .D(mem_rdata_latched_18_), .Q(mem_rdata_q_18_) );
DFFPOSX1 DFFPOSX1_979 ( .CLK(clk_bF_buf117), .D(mem_rdata_latched_19_), .Q(mem_rdata_q_19_) );
DFFPOSX1 DFFPOSX1_980 ( .CLK(clk_bF_buf116), .D(mem_rdata_latched_20_), .Q(mem_rdata_q_20_) );
DFFPOSX1 DFFPOSX1_981 ( .CLK(clk_bF_buf115), .D(mem_rdata_latched_21_), .Q(mem_rdata_q_21_) );
DFFPOSX1 DFFPOSX1_982 ( .CLK(clk_bF_buf114), .D(mem_rdata_latched_22_), .Q(mem_rdata_q_22_) );
DFFPOSX1 DFFPOSX1_983 ( .CLK(clk_bF_buf113), .D(mem_rdata_latched_23_), .Q(mem_rdata_q_23_) );
DFFPOSX1 DFFPOSX1_984 ( .CLK(clk_bF_buf112), .D(mem_rdata_latched_24_), .Q(mem_rdata_q_24_) );
DFFPOSX1 DFFPOSX1_985 ( .CLK(clk_bF_buf111), .D(mem_rdata_latched_25_), .Q(mem_rdata_q_25_) );
DFFPOSX1 DFFPOSX1_986 ( .CLK(clk_bF_buf110), .D(mem_rdata_latched_26_), .Q(mem_rdata_q_26_) );
DFFPOSX1 DFFPOSX1_987 ( .CLK(clk_bF_buf109), .D(mem_rdata_latched_27_), .Q(mem_rdata_q_27_) );
DFFPOSX1 DFFPOSX1_988 ( .CLK(clk_bF_buf108), .D(mem_rdata_latched_28_), .Q(mem_rdata_q_28_) );
DFFPOSX1 DFFPOSX1_989 ( .CLK(clk_bF_buf107), .D(mem_rdata_latched_29_), .Q(mem_rdata_q_29_) );
DFFPOSX1 DFFPOSX1_990 ( .CLK(clk_bF_buf106), .D(mem_rdata_latched_30_), .Q(mem_rdata_q_30_) );
DFFPOSX1 DFFPOSX1_991 ( .CLK(clk_bF_buf105), .D(mem_rdata_latched_31_), .Q(mem_rdata_q_31_) );
DFFPOSX1 DFFPOSX1_992 ( .CLK(clk_bF_buf104), .D(_6__0_), .Q(decoded_rs2_0_) );
DFFPOSX1 DFFPOSX1_993 ( .CLK(clk_bF_buf103), .D(_6__1_), .Q(decoded_rs2_1_) );
DFFPOSX1 DFFPOSX1_994 ( .CLK(clk_bF_buf102), .D(_6__2_), .Q(decoded_rs2_2_) );
DFFPOSX1 DFFPOSX1_995 ( .CLK(clk_bF_buf101), .D(_6__3_), .Q(decoded_rs2_3_) );
DFFPOSX1 DFFPOSX1_996 ( .CLK(clk_bF_buf100), .D(_6__4_), .Q(decoded_rs2_4_) );
DFFPOSX1 DFFPOSX1_997 ( .CLK(clk_bF_buf99), .D(_88_), .Q(cpu_state_0_) );
DFFPOSX1 DFFPOSX1_998 ( .CLK(clk_bF_buf98), .D(_93_), .Q(cpu_state_1_) );
DFFPOSX1 DFFPOSX1_999 ( .CLK(clk_bF_buf97), .D(_94_), .Q(cpu_state_2_) );
DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk_bF_buf96), .D(_89_), .Q(cpu_state_3_) );
DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk_bF_buf95), .D(_90_), .Q(cpu_state_4_) );
DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk_bF_buf94), .D(_91_), .Q(cpu_state_5_) );
DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk_bF_buf93), .D(_92_), .Q(cpu_state_6_) );
DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk_bF_buf92), .D(_1115_), .Q(cpuregs_8_[0]) );
DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk_bF_buf91), .D(_1116_), .Q(cpuregs_8_[1]) );
DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk_bF_buf90), .D(_1117_), .Q(cpuregs_8_[2]) );
DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk_bF_buf89), .D(_1118_), .Q(cpuregs_8_[3]) );
DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk_bF_buf88), .D(_1119_), .Q(cpuregs_8_[4]) );
DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk_bF_buf87), .D(_95_), .Q(cpuregs_8_[5]) );
DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk_bF_buf86), .D(_96_), .Q(cpuregs_8_[6]) );
DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk_bF_buf85), .D(_97_), .Q(cpuregs_8_[7]) );
DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk_bF_buf84), .D(_98_), .Q(cpuregs_8_[8]) );
DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk_bF_buf83), .D(_99_), .Q(cpuregs_8_[9]) );
DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk_bF_buf82), .D(_100_), .Q(cpuregs_8_[10]) );
DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk_bF_buf81), .D(_101_), .Q(cpuregs_8_[11]) );
DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk_bF_buf80), .D(_102_), .Q(cpuregs_8_[12]) );
DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk_bF_buf79), .D(_103_), .Q(cpuregs_8_[13]) );
DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk_bF_buf78), .D(_104_), .Q(cpuregs_8_[14]) );
DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk_bF_buf77), .D(_105_), .Q(cpuregs_8_[15]) );
DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk_bF_buf76), .D(_106_), .Q(cpuregs_8_[16]) );
DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk_bF_buf75), .D(_107_), .Q(cpuregs_8_[17]) );
DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk_bF_buf74), .D(_108_), .Q(cpuregs_8_[18]) );
DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk_bF_buf73), .D(_109_), .Q(cpuregs_8_[19]) );
DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk_bF_buf72), .D(_110_), .Q(cpuregs_8_[20]) );
DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk_bF_buf71), .D(_111_), .Q(cpuregs_8_[21]) );
DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk_bF_buf70), .D(_112_), .Q(cpuregs_8_[22]) );
DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk_bF_buf69), .D(_113_), .Q(cpuregs_8_[23]) );
DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk_bF_buf68), .D(_114_), .Q(cpuregs_8_[24]) );
DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk_bF_buf67), .D(_115_), .Q(cpuregs_8_[25]) );
DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk_bF_buf66), .D(_116_), .Q(cpuregs_8_[26]) );
DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk_bF_buf65), .D(_117_), .Q(cpuregs_8_[27]) );
DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk_bF_buf64), .D(_118_), .Q(cpuregs_8_[28]) );
DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk_bF_buf63), .D(_119_), .Q(cpuregs_8_[29]) );
DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk_bF_buf62), .D(_120_), .Q(cpuregs_8_[30]) );
DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk_bF_buf61), .D(_121_), .Q(cpuregs_8_[31]) );
DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk_bF_buf60), .D(_699_), .Q(cpuregs_21_[0]) );
DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk_bF_buf59), .D(_700_), .Q(cpuregs_21_[1]) );
DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk_bF_buf58), .D(_701_), .Q(cpuregs_21_[2]) );
DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk_bF_buf57), .D(_702_), .Q(cpuregs_21_[3]) );
DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk_bF_buf56), .D(_703_), .Q(cpuregs_21_[4]) );
DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk_bF_buf55), .D(_704_), .Q(cpuregs_21_[5]) );
DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk_bF_buf54), .D(_705_), .Q(cpuregs_21_[6]) );
DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk_bF_buf53), .D(_706_), .Q(cpuregs_21_[7]) );
DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk_bF_buf52), .D(_707_), .Q(cpuregs_21_[8]) );
DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk_bF_buf51), .D(_708_), .Q(cpuregs_21_[9]) );
DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk_bF_buf50), .D(_709_), .Q(cpuregs_21_[10]) );
DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk_bF_buf49), .D(_710_), .Q(cpuregs_21_[11]) );
DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk_bF_buf48), .D(_711_), .Q(cpuregs_21_[12]) );
DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk_bF_buf47), .D(_712_), .Q(cpuregs_21_[13]) );
DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk_bF_buf46), .D(_713_), .Q(cpuregs_21_[14]) );
DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk_bF_buf45), .D(_714_), .Q(cpuregs_21_[15]) );
DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk_bF_buf44), .D(_715_), .Q(cpuregs_21_[16]) );
DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk_bF_buf43), .D(_716_), .Q(cpuregs_21_[17]) );
DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk_bF_buf42), .D(_717_), .Q(cpuregs_21_[18]) );
DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk_bF_buf41), .D(_718_), .Q(cpuregs_21_[19]) );
DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk_bF_buf40), .D(_719_), .Q(cpuregs_21_[20]) );
DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk_bF_buf39), .D(_720_), .Q(cpuregs_21_[21]) );
DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk_bF_buf38), .D(_721_), .Q(cpuregs_21_[22]) );
DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk_bF_buf37), .D(_722_), .Q(cpuregs_21_[23]) );
DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk_bF_buf36), .D(_723_), .Q(cpuregs_21_[24]) );
DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk_bF_buf35), .D(_724_), .Q(cpuregs_21_[25]) );
DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk_bF_buf34), .D(_725_), .Q(cpuregs_21_[26]) );
DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk_bF_buf33), .D(_726_), .Q(cpuregs_21_[27]) );
DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk_bF_buf32), .D(_727_), .Q(cpuregs_21_[28]) );
DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk_bF_buf31), .D(_728_), .Q(cpuregs_21_[29]) );
DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk_bF_buf30), .D(_729_), .Q(cpuregs_21_[30]) );
DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk_bF_buf29), .D(_730_), .Q(cpuregs_21_[31]) );
DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk_bF_buf28), .D(_475_), .Q(cpuregs_28_[0]) );
DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk_bF_buf27), .D(_476_), .Q(cpuregs_28_[1]) );
DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk_bF_buf26), .D(_477_), .Q(cpuregs_28_[2]) );
DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk_bF_buf25), .D(_478_), .Q(cpuregs_28_[3]) );
DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk_bF_buf24), .D(_479_), .Q(cpuregs_28_[4]) );
DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk_bF_buf23), .D(_480_), .Q(cpuregs_28_[5]) );
DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk_bF_buf22), .D(_481_), .Q(cpuregs_28_[6]) );
DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk_bF_buf21), .D(_482_), .Q(cpuregs_28_[7]) );
DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk_bF_buf20), .D(_483_), .Q(cpuregs_28_[8]) );
DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk_bF_buf19), .D(_484_), .Q(cpuregs_28_[9]) );
DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk_bF_buf18), .D(_485_), .Q(cpuregs_28_[10]) );
DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk_bF_buf17), .D(_486_), .Q(cpuregs_28_[11]) );
DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk_bF_buf16), .D(_487_), .Q(cpuregs_28_[12]) );
DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk_bF_buf15), .D(_488_), .Q(cpuregs_28_[13]) );
DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk_bF_buf14), .D(_489_), .Q(cpuregs_28_[14]) );
DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk_bF_buf13), .D(_490_), .Q(cpuregs_28_[15]) );
DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk_bF_buf12), .D(_491_), .Q(cpuregs_28_[16]) );
DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk_bF_buf11), .D(_492_), .Q(cpuregs_28_[17]) );
DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk_bF_buf10), .D(_493_), .Q(cpuregs_28_[18]) );
DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk_bF_buf9), .D(_494_), .Q(cpuregs_28_[19]) );
DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk_bF_buf8), .D(_495_), .Q(cpuregs_28_[20]) );
DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk_bF_buf7), .D(_496_), .Q(cpuregs_28_[21]) );
DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk_bF_buf6), .D(_497_), .Q(cpuregs_28_[22]) );
DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk_bF_buf5), .D(_498_), .Q(cpuregs_28_[23]) );
DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk_bF_buf4), .D(_499_), .Q(cpuregs_28_[24]) );
DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk_bF_buf3), .D(_500_), .Q(cpuregs_28_[25]) );
DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk_bF_buf2), .D(_501_), .Q(cpuregs_28_[26]) );
DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk_bF_buf1), .D(_502_), .Q(cpuregs_28_[27]) );
DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk_bF_buf0), .D(_503_), .Q(cpuregs_28_[28]) );
DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk_bF_buf136), .D(_504_), .Q(cpuregs_28_[29]) );
DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk_bF_buf135), .D(_505_), .Q(cpuregs_28_[30]) );
DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk_bF_buf134), .D(_506_), .Q(cpuregs_28_[31]) );
DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk_bF_buf133), .D(_346_), .Q(cpuregs_0_[0]) );
DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk_bF_buf132), .D(_347_), .Q(cpuregs_0_[1]) );
DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk_bF_buf131), .D(_348_), .Q(cpuregs_0_[2]) );
DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk_bF_buf130), .D(_349_), .Q(cpuregs_0_[3]) );
DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk_bF_buf129), .D(_350_), .Q(cpuregs_0_[4]) );
DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk_bF_buf128), .D(_351_), .Q(cpuregs_0_[5]) );
DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk_bF_buf127), .D(_352_), .Q(cpuregs_0_[6]) );
DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk_bF_buf126), .D(_353_), .Q(cpuregs_0_[7]) );
DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk_bF_buf125), .D(_354_), .Q(cpuregs_0_[8]) );
DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk_bF_buf124), .D(_355_), .Q(cpuregs_0_[9]) );
DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk_bF_buf123), .D(_356_), .Q(cpuregs_0_[10]) );
DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk_bF_buf122), .D(_357_), .Q(cpuregs_0_[11]) );
DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk_bF_buf121), .D(_358_), .Q(cpuregs_0_[12]) );
DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk_bF_buf120), .D(_359_), .Q(cpuregs_0_[13]) );
DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk_bF_buf119), .D(_360_), .Q(cpuregs_0_[14]) );
DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk_bF_buf118), .D(_361_), .Q(cpuregs_0_[15]) );
DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk_bF_buf117), .D(_362_), .Q(cpuregs_0_[16]) );
DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk_bF_buf116), .D(_363_), .Q(cpuregs_0_[17]) );
DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk_bF_buf115), .D(_364_), .Q(cpuregs_0_[18]) );
DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk_bF_buf114), .D(_365_), .Q(cpuregs_0_[19]) );
DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk_bF_buf113), .D(_366_), .Q(cpuregs_0_[20]) );
DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk_bF_buf112), .D(_367_), .Q(cpuregs_0_[21]) );
DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk_bF_buf111), .D(_368_), .Q(cpuregs_0_[22]) );
DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk_bF_buf110), .D(_369_), .Q(cpuregs_0_[23]) );
DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk_bF_buf109), .D(_370_), .Q(cpuregs_0_[24]) );
DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk_bF_buf108), .D(_371_), .Q(cpuregs_0_[25]) );
DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk_bF_buf107), .D(_372_), .Q(cpuregs_0_[26]) );
DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk_bF_buf106), .D(_373_), .Q(cpuregs_0_[27]) );
DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk_bF_buf105), .D(_374_), .Q(cpuregs_0_[28]) );
DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk_bF_buf104), .D(_375_), .Q(cpuregs_0_[29]) );
DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk_bF_buf103), .D(_376_), .Q(cpuregs_0_[30]) );
DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk_bF_buf102), .D(_377_), .Q(cpuregs_0_[31]) );
DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk_bF_buf101), .D(_987_), .Q(cpuregs_16_[0]) );
DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk_bF_buf100), .D(_988_), .Q(cpuregs_16_[1]) );
DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk_bF_buf99), .D(_989_), .Q(cpuregs_16_[2]) );
DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk_bF_buf98), .D(_990_), .Q(cpuregs_16_[3]) );
DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk_bF_buf97), .D(_991_), .Q(cpuregs_16_[4]) );
DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk_bF_buf96), .D(_992_), .Q(cpuregs_16_[5]) );
DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk_bF_buf95), .D(_993_), .Q(cpuregs_16_[6]) );
DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk_bF_buf94), .D(_994_), .Q(cpuregs_16_[7]) );
DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk_bF_buf93), .D(_995_), .Q(cpuregs_16_[8]) );
DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk_bF_buf92), .D(_996_), .Q(cpuregs_16_[9]) );
DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk_bF_buf91), .D(_997_), .Q(cpuregs_16_[10]) );
DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk_bF_buf90), .D(_998_), .Q(cpuregs_16_[11]) );
DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk_bF_buf89), .D(_999_), .Q(cpuregs_16_[12]) );
DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk_bF_buf88), .D(_1000_), .Q(cpuregs_16_[13]) );
DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk_bF_buf87), .D(_1001_), .Q(cpuregs_16_[14]) );
DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk_bF_buf86), .D(_1002_), .Q(cpuregs_16_[15]) );
DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk_bF_buf85), .D(_1003_), .Q(cpuregs_16_[16]) );
DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk_bF_buf84), .D(_1004_), .Q(cpuregs_16_[17]) );
DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk_bF_buf83), .D(_1005_), .Q(cpuregs_16_[18]) );
DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk_bF_buf82), .D(_1006_), .Q(cpuregs_16_[19]) );
DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk_bF_buf81), .D(_1007_), .Q(cpuregs_16_[20]) );
DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk_bF_buf80), .D(_1008_), .Q(cpuregs_16_[21]) );
DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk_bF_buf79), .D(_1009_), .Q(cpuregs_16_[22]) );
DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk_bF_buf78), .D(_1010_), .Q(cpuregs_16_[23]) );
DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk_bF_buf77), .D(_1011_), .Q(cpuregs_16_[24]) );
DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk_bF_buf76), .D(_1012_), .Q(cpuregs_16_[25]) );
DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk_bF_buf75), .D(_1013_), .Q(cpuregs_16_[26]) );
DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk_bF_buf74), .D(_1014_), .Q(cpuregs_16_[27]) );
DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk_bF_buf73), .D(_1015_), .Q(cpuregs_16_[28]) );
DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk_bF_buf72), .D(_1016_), .Q(cpuregs_16_[29]) );
DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk_bF_buf71), .D(_1017_), .Q(cpuregs_16_[30]) );
DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk_bF_buf70), .D(_1018_), .Q(cpuregs_16_[31]) );
DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk_bF_buf69), .D(_827_), .Q(cpuregs_20_[0]) );
DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk_bF_buf68), .D(_828_), .Q(cpuregs_20_[1]) );
DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk_bF_buf67), .D(_829_), .Q(cpuregs_20_[2]) );
DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk_bF_buf66), .D(_830_), .Q(cpuregs_20_[3]) );
DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk_bF_buf65), .D(_831_), .Q(cpuregs_20_[4]) );
DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk_bF_buf64), .D(_832_), .Q(cpuregs_20_[5]) );
DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk_bF_buf63), .D(_833_), .Q(cpuregs_20_[6]) );
DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk_bF_buf62), .D(_834_), .Q(cpuregs_20_[7]) );
DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk_bF_buf61), .D(_835_), .Q(cpuregs_20_[8]) );
DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk_bF_buf60), .D(_836_), .Q(cpuregs_20_[9]) );
DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk_bF_buf59), .D(_837_), .Q(cpuregs_20_[10]) );
DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk_bF_buf58), .D(_838_), .Q(cpuregs_20_[11]) );
DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk_bF_buf57), .D(_839_), .Q(cpuregs_20_[12]) );
DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk_bF_buf56), .D(_840_), .Q(cpuregs_20_[13]) );
DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk_bF_buf55), .D(_841_), .Q(cpuregs_20_[14]) );
DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk_bF_buf54), .D(_842_), .Q(cpuregs_20_[15]) );
DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk_bF_buf53), .D(_843_), .Q(cpuregs_20_[16]) );
DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk_bF_buf52), .D(_844_), .Q(cpuregs_20_[17]) );
DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk_bF_buf51), .D(_845_), .Q(cpuregs_20_[18]) );
DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk_bF_buf50), .D(_846_), .Q(cpuregs_20_[19]) );
DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk_bF_buf49), .D(_847_), .Q(cpuregs_20_[20]) );
DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk_bF_buf48), .D(_848_), .Q(cpuregs_20_[21]) );
DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk_bF_buf47), .D(_849_), .Q(cpuregs_20_[22]) );
DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk_bF_buf46), .D(_850_), .Q(cpuregs_20_[23]) );
DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk_bF_buf45), .D(_851_), .Q(cpuregs_20_[24]) );
DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk_bF_buf44), .D(_852_), .Q(cpuregs_20_[25]) );
DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk_bF_buf43), .D(_853_), .Q(cpuregs_20_[26]) );
DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk_bF_buf42), .D(_854_), .Q(cpuregs_20_[27]) );
DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk_bF_buf41), .D(_855_), .Q(cpuregs_20_[28]) );
DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk_bF_buf40), .D(_856_), .Q(cpuregs_20_[29]) );
DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk_bF_buf39), .D(_857_), .Q(cpuregs_20_[30]) );
DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk_bF_buf38), .D(_858_), .Q(cpuregs_20_[31]) );
DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk_bF_buf37), .D(_507_), .Q(cpuregs_27_[0]) );
DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk_bF_buf36), .D(_508_), .Q(cpuregs_27_[1]) );
DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk_bF_buf35), .D(_509_), .Q(cpuregs_27_[2]) );
DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk_bF_buf34), .D(_510_), .Q(cpuregs_27_[3]) );
DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk_bF_buf33), .D(_511_), .Q(cpuregs_27_[4]) );
DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk_bF_buf32), .D(_512_), .Q(cpuregs_27_[5]) );
DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk_bF_buf31), .D(_513_), .Q(cpuregs_27_[6]) );
DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk_bF_buf30), .D(_514_), .Q(cpuregs_27_[7]) );
DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk_bF_buf29), .D(_515_), .Q(cpuregs_27_[8]) );
DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk_bF_buf28), .D(_516_), .Q(cpuregs_27_[9]) );
DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk_bF_buf27), .D(_517_), .Q(cpuregs_27_[10]) );
DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk_bF_buf26), .D(_518_), .Q(cpuregs_27_[11]) );
DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk_bF_buf25), .D(_519_), .Q(cpuregs_27_[12]) );
DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk_bF_buf24), .D(_520_), .Q(cpuregs_27_[13]) );
DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk_bF_buf23), .D(_521_), .Q(cpuregs_27_[14]) );
DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk_bF_buf22), .D(_522_), .Q(cpuregs_27_[15]) );
DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk_bF_buf21), .D(_523_), .Q(cpuregs_27_[16]) );
DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk_bF_buf20), .D(_524_), .Q(cpuregs_27_[17]) );
DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk_bF_buf19), .D(_525_), .Q(cpuregs_27_[18]) );
DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk_bF_buf18), .D(_526_), .Q(cpuregs_27_[19]) );
DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk_bF_buf17), .D(_527_), .Q(cpuregs_27_[20]) );
DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk_bF_buf16), .D(_528_), .Q(cpuregs_27_[21]) );
DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk_bF_buf15), .D(_529_), .Q(cpuregs_27_[22]) );
DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk_bF_buf14), .D(_530_), .Q(cpuregs_27_[23]) );
DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk_bF_buf13), .D(_531_), .Q(cpuregs_27_[24]) );
DFFPOSX1 DFFPOSX1_1221 ( .CLK(clk_bF_buf12), .D(_532_), .Q(cpuregs_27_[25]) );
DFFPOSX1 DFFPOSX1_1222 ( .CLK(clk_bF_buf11), .D(_533_), .Q(cpuregs_27_[26]) );
DFFPOSX1 DFFPOSX1_1223 ( .CLK(clk_bF_buf10), .D(_534_), .Q(cpuregs_27_[27]) );
DFFPOSX1 DFFPOSX1_1224 ( .CLK(clk_bF_buf9), .D(_535_), .Q(cpuregs_27_[28]) );
DFFPOSX1 DFFPOSX1_1225 ( .CLK(clk_bF_buf8), .D(_536_), .Q(cpuregs_27_[29]) );
DFFPOSX1 DFFPOSX1_1226 ( .CLK(clk_bF_buf7), .D(_537_), .Q(cpuregs_27_[30]) );
DFFPOSX1 DFFPOSX1_1227 ( .CLK(clk_bF_buf6), .D(_538_), .Q(cpuregs_27_[31]) );
DFFPOSX1 DFFPOSX1_1228 ( .CLK(clk_bF_buf5), .D(_443_), .Q(cpuregs_29_[0]) );
DFFPOSX1 DFFPOSX1_1229 ( .CLK(clk_bF_buf4), .D(_444_), .Q(cpuregs_29_[1]) );
DFFPOSX1 DFFPOSX1_1230 ( .CLK(clk_bF_buf3), .D(_445_), .Q(cpuregs_29_[2]) );
DFFPOSX1 DFFPOSX1_1231 ( .CLK(clk_bF_buf2), .D(_446_), .Q(cpuregs_29_[3]) );
DFFPOSX1 DFFPOSX1_1232 ( .CLK(clk_bF_buf1), .D(_447_), .Q(cpuregs_29_[4]) );
DFFPOSX1 DFFPOSX1_1233 ( .CLK(clk_bF_buf0), .D(_448_), .Q(cpuregs_29_[5]) );
DFFPOSX1 DFFPOSX1_1234 ( .CLK(clk_bF_buf136), .D(_449_), .Q(cpuregs_29_[6]) );
DFFPOSX1 DFFPOSX1_1235 ( .CLK(clk_bF_buf135), .D(_450_), .Q(cpuregs_29_[7]) );
DFFPOSX1 DFFPOSX1_1236 ( .CLK(clk_bF_buf134), .D(_451_), .Q(cpuregs_29_[8]) );
DFFPOSX1 DFFPOSX1_1237 ( .CLK(clk_bF_buf133), .D(_452_), .Q(cpuregs_29_[9]) );
DFFPOSX1 DFFPOSX1_1238 ( .CLK(clk_bF_buf132), .D(_453_), .Q(cpuregs_29_[10]) );
DFFPOSX1 DFFPOSX1_1239 ( .CLK(clk_bF_buf131), .D(_454_), .Q(cpuregs_29_[11]) );
DFFPOSX1 DFFPOSX1_1240 ( .CLK(clk_bF_buf130), .D(_455_), .Q(cpuregs_29_[12]) );
DFFPOSX1 DFFPOSX1_1241 ( .CLK(clk_bF_buf129), .D(_456_), .Q(cpuregs_29_[13]) );
DFFPOSX1 DFFPOSX1_1242 ( .CLK(clk_bF_buf128), .D(_457_), .Q(cpuregs_29_[14]) );
DFFPOSX1 DFFPOSX1_1243 ( .CLK(clk_bF_buf127), .D(_458_), .Q(cpuregs_29_[15]) );
DFFPOSX1 DFFPOSX1_1244 ( .CLK(clk_bF_buf126), .D(_459_), .Q(cpuregs_29_[16]) );
DFFPOSX1 DFFPOSX1_1245 ( .CLK(clk_bF_buf125), .D(_460_), .Q(cpuregs_29_[17]) );
DFFPOSX1 DFFPOSX1_1246 ( .CLK(clk_bF_buf124), .D(_461_), .Q(cpuregs_29_[18]) );
DFFPOSX1 DFFPOSX1_1247 ( .CLK(clk_bF_buf123), .D(_462_), .Q(cpuregs_29_[19]) );
DFFPOSX1 DFFPOSX1_1248 ( .CLK(clk_bF_buf122), .D(_463_), .Q(cpuregs_29_[20]) );
DFFPOSX1 DFFPOSX1_1249 ( .CLK(clk_bF_buf121), .D(_464_), .Q(cpuregs_29_[21]) );
DFFPOSX1 DFFPOSX1_1250 ( .CLK(clk_bF_buf120), .D(_465_), .Q(cpuregs_29_[22]) );
DFFPOSX1 DFFPOSX1_1251 ( .CLK(clk_bF_buf119), .D(_466_), .Q(cpuregs_29_[23]) );
DFFPOSX1 DFFPOSX1_1252 ( .CLK(clk_bF_buf118), .D(_467_), .Q(cpuregs_29_[24]) );
DFFPOSX1 DFFPOSX1_1253 ( .CLK(clk_bF_buf117), .D(_468_), .Q(cpuregs_29_[25]) );
DFFPOSX1 DFFPOSX1_1254 ( .CLK(clk_bF_buf116), .D(_469_), .Q(cpuregs_29_[26]) );
DFFPOSX1 DFFPOSX1_1255 ( .CLK(clk_bF_buf115), .D(_470_), .Q(cpuregs_29_[27]) );
DFFPOSX1 DFFPOSX1_1256 ( .CLK(clk_bF_buf114), .D(_471_), .Q(cpuregs_29_[28]) );
DFFPOSX1 DFFPOSX1_1257 ( .CLK(clk_bF_buf113), .D(_472_), .Q(cpuregs_29_[29]) );
DFFPOSX1 DFFPOSX1_1258 ( .CLK(clk_bF_buf112), .D(_473_), .Q(cpuregs_29_[30]) );
DFFPOSX1 DFFPOSX1_1259 ( .CLK(clk_bF_buf111), .D(_474_), .Q(cpuregs_29_[31]) );
DFFPOSX1 DFFPOSX1_1260 ( .CLK(clk_bF_buf110), .D(_1019_), .Q(cpuregs_15_[0]) );
DFFPOSX1 DFFPOSX1_1261 ( .CLK(clk_bF_buf109), .D(_1020_), .Q(cpuregs_15_[1]) );
DFFPOSX1 DFFPOSX1_1262 ( .CLK(clk_bF_buf108), .D(_1021_), .Q(cpuregs_15_[2]) );
DFFPOSX1 DFFPOSX1_1263 ( .CLK(clk_bF_buf107), .D(_1022_), .Q(cpuregs_15_[3]) );
DFFPOSX1 DFFPOSX1_1264 ( .CLK(clk_bF_buf106), .D(_1023_), .Q(cpuregs_15_[4]) );
DFFPOSX1 DFFPOSX1_1265 ( .CLK(clk_bF_buf105), .D(_1024_), .Q(cpuregs_15_[5]) );
DFFPOSX1 DFFPOSX1_1266 ( .CLK(clk_bF_buf104), .D(_1025_), .Q(cpuregs_15_[6]) );
DFFPOSX1 DFFPOSX1_1267 ( .CLK(clk_bF_buf103), .D(_1026_), .Q(cpuregs_15_[7]) );
DFFPOSX1 DFFPOSX1_1268 ( .CLK(clk_bF_buf102), .D(_1027_), .Q(cpuregs_15_[8]) );
DFFPOSX1 DFFPOSX1_1269 ( .CLK(clk_bF_buf101), .D(_1028_), .Q(cpuregs_15_[9]) );
DFFPOSX1 DFFPOSX1_1270 ( .CLK(clk_bF_buf100), .D(_1029_), .Q(cpuregs_15_[10]) );
DFFPOSX1 DFFPOSX1_1271 ( .CLK(clk_bF_buf99), .D(_1030_), .Q(cpuregs_15_[11]) );
DFFPOSX1 DFFPOSX1_1272 ( .CLK(clk_bF_buf98), .D(_1031_), .Q(cpuregs_15_[12]) );
DFFPOSX1 DFFPOSX1_1273 ( .CLK(clk_bF_buf97), .D(_1032_), .Q(cpuregs_15_[13]) );
DFFPOSX1 DFFPOSX1_1274 ( .CLK(clk_bF_buf96), .D(_1033_), .Q(cpuregs_15_[14]) );
DFFPOSX1 DFFPOSX1_1275 ( .CLK(clk_bF_buf95), .D(_1034_), .Q(cpuregs_15_[15]) );
DFFPOSX1 DFFPOSX1_1276 ( .CLK(clk_bF_buf94), .D(_1035_), .Q(cpuregs_15_[16]) );
DFFPOSX1 DFFPOSX1_1277 ( .CLK(clk_bF_buf93), .D(_1036_), .Q(cpuregs_15_[17]) );
DFFPOSX1 DFFPOSX1_1278 ( .CLK(clk_bF_buf92), .D(_1037_), .Q(cpuregs_15_[18]) );
DFFPOSX1 DFFPOSX1_1279 ( .CLK(clk_bF_buf91), .D(_1038_), .Q(cpuregs_15_[19]) );
DFFPOSX1 DFFPOSX1_1280 ( .CLK(clk_bF_buf90), .D(_1039_), .Q(cpuregs_15_[20]) );
DFFPOSX1 DFFPOSX1_1281 ( .CLK(clk_bF_buf89), .D(_1040_), .Q(cpuregs_15_[21]) );
DFFPOSX1 DFFPOSX1_1282 ( .CLK(clk_bF_buf88), .D(_1041_), .Q(cpuregs_15_[22]) );
DFFPOSX1 DFFPOSX1_1283 ( .CLK(clk_bF_buf87), .D(_1042_), .Q(cpuregs_15_[23]) );
DFFPOSX1 DFFPOSX1_1284 ( .CLK(clk_bF_buf86), .D(_1043_), .Q(cpuregs_15_[24]) );
DFFPOSX1 DFFPOSX1_1285 ( .CLK(clk_bF_buf85), .D(_1044_), .Q(cpuregs_15_[25]) );
DFFPOSX1 DFFPOSX1_1286 ( .CLK(clk_bF_buf84), .D(_1045_), .Q(cpuregs_15_[26]) );
DFFPOSX1 DFFPOSX1_1287 ( .CLK(clk_bF_buf83), .D(_1046_), .Q(cpuregs_15_[27]) );
DFFPOSX1 DFFPOSX1_1288 ( .CLK(clk_bF_buf82), .D(_1047_), .Q(cpuregs_15_[28]) );
DFFPOSX1 DFFPOSX1_1289 ( .CLK(clk_bF_buf81), .D(_1048_), .Q(cpuregs_15_[29]) );
DFFPOSX1 DFFPOSX1_1290 ( .CLK(clk_bF_buf80), .D(_1049_), .Q(cpuregs_15_[30]) );
DFFPOSX1 DFFPOSX1_1291 ( .CLK(clk_bF_buf79), .D(_1050_), .Q(cpuregs_15_[31]) );
DFFPOSX1 DFFPOSX1_1292 ( .CLK(clk_bF_buf78), .D(_1051_), .Q(cpuregs_14_[0]) );
DFFPOSX1 DFFPOSX1_1293 ( .CLK(clk_bF_buf77), .D(_1052_), .Q(cpuregs_14_[1]) );
DFFPOSX1 DFFPOSX1_1294 ( .CLK(clk_bF_buf76), .D(_1053_), .Q(cpuregs_14_[2]) );
DFFPOSX1 DFFPOSX1_1295 ( .CLK(clk_bF_buf75), .D(_1054_), .Q(cpuregs_14_[3]) );
DFFPOSX1 DFFPOSX1_1296 ( .CLK(clk_bF_buf74), .D(_1055_), .Q(cpuregs_14_[4]) );
DFFPOSX1 DFFPOSX1_1297 ( .CLK(clk_bF_buf73), .D(_1056_), .Q(cpuregs_14_[5]) );
DFFPOSX1 DFFPOSX1_1298 ( .CLK(clk_bF_buf72), .D(_1057_), .Q(cpuregs_14_[6]) );
DFFPOSX1 DFFPOSX1_1299 ( .CLK(clk_bF_buf71), .D(_1058_), .Q(cpuregs_14_[7]) );
DFFPOSX1 DFFPOSX1_1300 ( .CLK(clk_bF_buf70), .D(_1059_), .Q(cpuregs_14_[8]) );
DFFPOSX1 DFFPOSX1_1301 ( .CLK(clk_bF_buf69), .D(_1060_), .Q(cpuregs_14_[9]) );
DFFPOSX1 DFFPOSX1_1302 ( .CLK(clk_bF_buf68), .D(_1061_), .Q(cpuregs_14_[10]) );
DFFPOSX1 DFFPOSX1_1303 ( .CLK(clk_bF_buf67), .D(_1062_), .Q(cpuregs_14_[11]) );
DFFPOSX1 DFFPOSX1_1304 ( .CLK(clk_bF_buf66), .D(_1063_), .Q(cpuregs_14_[12]) );
DFFPOSX1 DFFPOSX1_1305 ( .CLK(clk_bF_buf65), .D(_1064_), .Q(cpuregs_14_[13]) );
DFFPOSX1 DFFPOSX1_1306 ( .CLK(clk_bF_buf64), .D(_1065_), .Q(cpuregs_14_[14]) );
DFFPOSX1 DFFPOSX1_1307 ( .CLK(clk_bF_buf63), .D(_1066_), .Q(cpuregs_14_[15]) );
DFFPOSX1 DFFPOSX1_1308 ( .CLK(clk_bF_buf62), .D(_1067_), .Q(cpuregs_14_[16]) );
DFFPOSX1 DFFPOSX1_1309 ( .CLK(clk_bF_buf61), .D(_1068_), .Q(cpuregs_14_[17]) );
DFFPOSX1 DFFPOSX1_1310 ( .CLK(clk_bF_buf60), .D(_1069_), .Q(cpuregs_14_[18]) );
DFFPOSX1 DFFPOSX1_1311 ( .CLK(clk_bF_buf59), .D(_1070_), .Q(cpuregs_14_[19]) );
DFFPOSX1 DFFPOSX1_1312 ( .CLK(clk_bF_buf58), .D(_1071_), .Q(cpuregs_14_[20]) );
DFFPOSX1 DFFPOSX1_1313 ( .CLK(clk_bF_buf57), .D(_1072_), .Q(cpuregs_14_[21]) );
DFFPOSX1 DFFPOSX1_1314 ( .CLK(clk_bF_buf56), .D(_1073_), .Q(cpuregs_14_[22]) );
DFFPOSX1 DFFPOSX1_1315 ( .CLK(clk_bF_buf55), .D(_1074_), .Q(cpuregs_14_[23]) );
DFFPOSX1 DFFPOSX1_1316 ( .CLK(clk_bF_buf54), .D(_1075_), .Q(cpuregs_14_[24]) );
DFFPOSX1 DFFPOSX1_1317 ( .CLK(clk_bF_buf53), .D(_1076_), .Q(cpuregs_14_[25]) );
DFFPOSX1 DFFPOSX1_1318 ( .CLK(clk_bF_buf52), .D(_1077_), .Q(cpuregs_14_[26]) );
DFFPOSX1 DFFPOSX1_1319 ( .CLK(clk_bF_buf51), .D(_1078_), .Q(cpuregs_14_[27]) );
DFFPOSX1 DFFPOSX1_1320 ( .CLK(clk_bF_buf50), .D(_1079_), .Q(cpuregs_14_[28]) );
DFFPOSX1 DFFPOSX1_1321 ( .CLK(clk_bF_buf49), .D(_1080_), .Q(cpuregs_14_[29]) );
DFFPOSX1 DFFPOSX1_1322 ( .CLK(clk_bF_buf48), .D(_1081_), .Q(cpuregs_14_[30]) );
DFFPOSX1 DFFPOSX1_1323 ( .CLK(clk_bF_buf47), .D(_1082_), .Q(cpuregs_14_[31]) );
DFFPOSX1 DFFPOSX1_1324 ( .CLK(clk_bF_buf46), .D(_955_), .Q(cpuregs_17_[0]) );
DFFPOSX1 DFFPOSX1_1325 ( .CLK(clk_bF_buf45), .D(_956_), .Q(cpuregs_17_[1]) );
DFFPOSX1 DFFPOSX1_1326 ( .CLK(clk_bF_buf44), .D(_957_), .Q(cpuregs_17_[2]) );
DFFPOSX1 DFFPOSX1_1327 ( .CLK(clk_bF_buf43), .D(_958_), .Q(cpuregs_17_[3]) );
DFFPOSX1 DFFPOSX1_1328 ( .CLK(clk_bF_buf42), .D(_959_), .Q(cpuregs_17_[4]) );
DFFPOSX1 DFFPOSX1_1329 ( .CLK(clk_bF_buf41), .D(_960_), .Q(cpuregs_17_[5]) );
DFFPOSX1 DFFPOSX1_1330 ( .CLK(clk_bF_buf40), .D(_961_), .Q(cpuregs_17_[6]) );
DFFPOSX1 DFFPOSX1_1331 ( .CLK(clk_bF_buf39), .D(_962_), .Q(cpuregs_17_[7]) );
DFFPOSX1 DFFPOSX1_1332 ( .CLK(clk_bF_buf38), .D(_963_), .Q(cpuregs_17_[8]) );
DFFPOSX1 DFFPOSX1_1333 ( .CLK(clk_bF_buf37), .D(_964_), .Q(cpuregs_17_[9]) );
DFFPOSX1 DFFPOSX1_1334 ( .CLK(clk_bF_buf36), .D(_965_), .Q(cpuregs_17_[10]) );
DFFPOSX1 DFFPOSX1_1335 ( .CLK(clk_bF_buf35), .D(_966_), .Q(cpuregs_17_[11]) );
DFFPOSX1 DFFPOSX1_1336 ( .CLK(clk_bF_buf34), .D(_967_), .Q(cpuregs_17_[12]) );
DFFPOSX1 DFFPOSX1_1337 ( .CLK(clk_bF_buf33), .D(_968_), .Q(cpuregs_17_[13]) );
DFFPOSX1 DFFPOSX1_1338 ( .CLK(clk_bF_buf32), .D(_969_), .Q(cpuregs_17_[14]) );
DFFPOSX1 DFFPOSX1_1339 ( .CLK(clk_bF_buf31), .D(_970_), .Q(cpuregs_17_[15]) );
DFFPOSX1 DFFPOSX1_1340 ( .CLK(clk_bF_buf30), .D(_971_), .Q(cpuregs_17_[16]) );
DFFPOSX1 DFFPOSX1_1341 ( .CLK(clk_bF_buf29), .D(_972_), .Q(cpuregs_17_[17]) );
DFFPOSX1 DFFPOSX1_1342 ( .CLK(clk_bF_buf28), .D(_973_), .Q(cpuregs_17_[18]) );
DFFPOSX1 DFFPOSX1_1343 ( .CLK(clk_bF_buf27), .D(_974_), .Q(cpuregs_17_[19]) );
DFFPOSX1 DFFPOSX1_1344 ( .CLK(clk_bF_buf26), .D(_975_), .Q(cpuregs_17_[20]) );
DFFPOSX1 DFFPOSX1_1345 ( .CLK(clk_bF_buf25), .D(_976_), .Q(cpuregs_17_[21]) );
DFFPOSX1 DFFPOSX1_1346 ( .CLK(clk_bF_buf24), .D(_977_), .Q(cpuregs_17_[22]) );
DFFPOSX1 DFFPOSX1_1347 ( .CLK(clk_bF_buf23), .D(_978_), .Q(cpuregs_17_[23]) );
DFFPOSX1 DFFPOSX1_1348 ( .CLK(clk_bF_buf22), .D(_979_), .Q(cpuregs_17_[24]) );
DFFPOSX1 DFFPOSX1_1349 ( .CLK(clk_bF_buf21), .D(_980_), .Q(cpuregs_17_[25]) );
DFFPOSX1 DFFPOSX1_1350 ( .CLK(clk_bF_buf20), .D(_981_), .Q(cpuregs_17_[26]) );
DFFPOSX1 DFFPOSX1_1351 ( .CLK(clk_bF_buf19), .D(_982_), .Q(cpuregs_17_[27]) );
DFFPOSX1 DFFPOSX1_1352 ( .CLK(clk_bF_buf18), .D(_983_), .Q(cpuregs_17_[28]) );
DFFPOSX1 DFFPOSX1_1353 ( .CLK(clk_bF_buf17), .D(_984_), .Q(cpuregs_17_[29]) );
DFFPOSX1 DFFPOSX1_1354 ( .CLK(clk_bF_buf16), .D(_985_), .Q(cpuregs_17_[30]) );
DFFPOSX1 DFFPOSX1_1355 ( .CLK(clk_bF_buf15), .D(_986_), .Q(cpuregs_17_[31]) );
DFFPOSX1 DFFPOSX1_1356 ( .CLK(clk_bF_buf14), .D(_314_), .Q(cpuregs_1_[0]) );
DFFPOSX1 DFFPOSX1_1357 ( .CLK(clk_bF_buf13), .D(_315_), .Q(cpuregs_1_[1]) );
DFFPOSX1 DFFPOSX1_1358 ( .CLK(clk_bF_buf12), .D(_316_), .Q(cpuregs_1_[2]) );
DFFPOSX1 DFFPOSX1_1359 ( .CLK(clk_bF_buf11), .D(_317_), .Q(cpuregs_1_[3]) );
DFFPOSX1 DFFPOSX1_1360 ( .CLK(clk_bF_buf10), .D(_318_), .Q(cpuregs_1_[4]) );
DFFPOSX1 DFFPOSX1_1361 ( .CLK(clk_bF_buf9), .D(_319_), .Q(cpuregs_1_[5]) );
DFFPOSX1 DFFPOSX1_1362 ( .CLK(clk_bF_buf8), .D(_320_), .Q(cpuregs_1_[6]) );
DFFPOSX1 DFFPOSX1_1363 ( .CLK(clk_bF_buf7), .D(_321_), .Q(cpuregs_1_[7]) );
DFFPOSX1 DFFPOSX1_1364 ( .CLK(clk_bF_buf6), .D(_322_), .Q(cpuregs_1_[8]) );
DFFPOSX1 DFFPOSX1_1365 ( .CLK(clk_bF_buf5), .D(_323_), .Q(cpuregs_1_[9]) );
DFFPOSX1 DFFPOSX1_1366 ( .CLK(clk_bF_buf4), .D(_324_), .Q(cpuregs_1_[10]) );
DFFPOSX1 DFFPOSX1_1367 ( .CLK(clk_bF_buf3), .D(_325_), .Q(cpuregs_1_[11]) );
DFFPOSX1 DFFPOSX1_1368 ( .CLK(clk_bF_buf2), .D(_326_), .Q(cpuregs_1_[12]) );
DFFPOSX1 DFFPOSX1_1369 ( .CLK(clk_bF_buf1), .D(_327_), .Q(cpuregs_1_[13]) );
DFFPOSX1 DFFPOSX1_1370 ( .CLK(clk_bF_buf0), .D(_328_), .Q(cpuregs_1_[14]) );
DFFPOSX1 DFFPOSX1_1371 ( .CLK(clk_bF_buf136), .D(_329_), .Q(cpuregs_1_[15]) );
DFFPOSX1 DFFPOSX1_1372 ( .CLK(clk_bF_buf135), .D(_330_), .Q(cpuregs_1_[16]) );
DFFPOSX1 DFFPOSX1_1373 ( .CLK(clk_bF_buf134), .D(_331_), .Q(cpuregs_1_[17]) );
DFFPOSX1 DFFPOSX1_1374 ( .CLK(clk_bF_buf133), .D(_332_), .Q(cpuregs_1_[18]) );
DFFPOSX1 DFFPOSX1_1375 ( .CLK(clk_bF_buf132), .D(_333_), .Q(cpuregs_1_[19]) );
DFFPOSX1 DFFPOSX1_1376 ( .CLK(clk_bF_buf131), .D(_334_), .Q(cpuregs_1_[20]) );
DFFPOSX1 DFFPOSX1_1377 ( .CLK(clk_bF_buf130), .D(_335_), .Q(cpuregs_1_[21]) );
DFFPOSX1 DFFPOSX1_1378 ( .CLK(clk_bF_buf129), .D(_336_), .Q(cpuregs_1_[22]) );
DFFPOSX1 DFFPOSX1_1379 ( .CLK(clk_bF_buf128), .D(_337_), .Q(cpuregs_1_[23]) );
DFFPOSX1 DFFPOSX1_1380 ( .CLK(clk_bF_buf127), .D(_338_), .Q(cpuregs_1_[24]) );
DFFPOSX1 DFFPOSX1_1381 ( .CLK(clk_bF_buf126), .D(_339_), .Q(cpuregs_1_[25]) );
DFFPOSX1 DFFPOSX1_1382 ( .CLK(clk_bF_buf125), .D(_340_), .Q(cpuregs_1_[26]) );
DFFPOSX1 DFFPOSX1_1383 ( .CLK(clk_bF_buf124), .D(_341_), .Q(cpuregs_1_[27]) );
DFFPOSX1 DFFPOSX1_1384 ( .CLK(clk_bF_buf123), .D(_342_), .Q(cpuregs_1_[28]) );
DFFPOSX1 DFFPOSX1_1385 ( .CLK(clk_bF_buf122), .D(_343_), .Q(cpuregs_1_[29]) );
DFFPOSX1 DFFPOSX1_1386 ( .CLK(clk_bF_buf121), .D(_344_), .Q(cpuregs_1_[30]) );
DFFPOSX1 DFFPOSX1_1387 ( .CLK(clk_bF_buf120), .D(_345_), .Q(cpuregs_1_[31]) );
DFFPOSX1 DFFPOSX1_1388 ( .CLK(clk_bF_buf119), .D(_378_), .Q(mem_wordsize_0_) );
DFFPOSX1 DFFPOSX1_1389 ( .CLK(clk_bF_buf118), .D(_87_), .Q(mem_wordsize_2_) );
DFFPOSX1 DFFPOSX1_1390 ( .CLK(clk_bF_buf117), .D(_923_), .Q(cpuregs_18_[0]) );
DFFPOSX1 DFFPOSX1_1391 ( .CLK(clk_bF_buf116), .D(_924_), .Q(cpuregs_18_[1]) );
DFFPOSX1 DFFPOSX1_1392 ( .CLK(clk_bF_buf115), .D(_925_), .Q(cpuregs_18_[2]) );
DFFPOSX1 DFFPOSX1_1393 ( .CLK(clk_bF_buf114), .D(_926_), .Q(cpuregs_18_[3]) );
DFFPOSX1 DFFPOSX1_1394 ( .CLK(clk_bF_buf113), .D(_927_), .Q(cpuregs_18_[4]) );
DFFPOSX1 DFFPOSX1_1395 ( .CLK(clk_bF_buf112), .D(_928_), .Q(cpuregs_18_[5]) );
DFFPOSX1 DFFPOSX1_1396 ( .CLK(clk_bF_buf111), .D(_929_), .Q(cpuregs_18_[6]) );
DFFPOSX1 DFFPOSX1_1397 ( .CLK(clk_bF_buf110), .D(_930_), .Q(cpuregs_18_[7]) );
DFFPOSX1 DFFPOSX1_1398 ( .CLK(clk_bF_buf109), .D(_931_), .Q(cpuregs_18_[8]) );
DFFPOSX1 DFFPOSX1_1399 ( .CLK(clk_bF_buf108), .D(_932_), .Q(cpuregs_18_[9]) );
DFFPOSX1 DFFPOSX1_1400 ( .CLK(clk_bF_buf107), .D(_933_), .Q(cpuregs_18_[10]) );
DFFPOSX1 DFFPOSX1_1401 ( .CLK(clk_bF_buf106), .D(_934_), .Q(cpuregs_18_[11]) );
DFFPOSX1 DFFPOSX1_1402 ( .CLK(clk_bF_buf105), .D(_935_), .Q(cpuregs_18_[12]) );
DFFPOSX1 DFFPOSX1_1403 ( .CLK(clk_bF_buf104), .D(_936_), .Q(cpuregs_18_[13]) );
DFFPOSX1 DFFPOSX1_1404 ( .CLK(clk_bF_buf103), .D(_937_), .Q(cpuregs_18_[14]) );
DFFPOSX1 DFFPOSX1_1405 ( .CLK(clk_bF_buf102), .D(_938_), .Q(cpuregs_18_[15]) );
DFFPOSX1 DFFPOSX1_1406 ( .CLK(clk_bF_buf101), .D(_939_), .Q(cpuregs_18_[16]) );
DFFPOSX1 DFFPOSX1_1407 ( .CLK(clk_bF_buf100), .D(_940_), .Q(cpuregs_18_[17]) );
DFFPOSX1 DFFPOSX1_1408 ( .CLK(clk_bF_buf99), .D(_941_), .Q(cpuregs_18_[18]) );
DFFPOSX1 DFFPOSX1_1409 ( .CLK(clk_bF_buf98), .D(_942_), .Q(cpuregs_18_[19]) );
DFFPOSX1 DFFPOSX1_1410 ( .CLK(clk_bF_buf97), .D(_943_), .Q(cpuregs_18_[20]) );
DFFPOSX1 DFFPOSX1_1411 ( .CLK(clk_bF_buf96), .D(_944_), .Q(cpuregs_18_[21]) );
DFFPOSX1 DFFPOSX1_1412 ( .CLK(clk_bF_buf95), .D(_945_), .Q(cpuregs_18_[22]) );
DFFPOSX1 DFFPOSX1_1413 ( .CLK(clk_bF_buf94), .D(_946_), .Q(cpuregs_18_[23]) );
DFFPOSX1 DFFPOSX1_1414 ( .CLK(clk_bF_buf93), .D(_947_), .Q(cpuregs_18_[24]) );
DFFPOSX1 DFFPOSX1_1415 ( .CLK(clk_bF_buf92), .D(_948_), .Q(cpuregs_18_[25]) );
DFFPOSX1 DFFPOSX1_1416 ( .CLK(clk_bF_buf91), .D(_949_), .Q(cpuregs_18_[26]) );
DFFPOSX1 DFFPOSX1_1417 ( .CLK(clk_bF_buf90), .D(_950_), .Q(cpuregs_18_[27]) );
DFFPOSX1 DFFPOSX1_1418 ( .CLK(clk_bF_buf89), .D(_951_), .Q(cpuregs_18_[28]) );
DFFPOSX1 DFFPOSX1_1419 ( .CLK(clk_bF_buf88), .D(_952_), .Q(cpuregs_18_[29]) );
DFFPOSX1 DFFPOSX1_1420 ( .CLK(clk_bF_buf87), .D(_953_), .Q(cpuregs_18_[30]) );
DFFPOSX1 DFFPOSX1_1421 ( .CLK(clk_bF_buf86), .D(_954_), .Q(cpuregs_18_[31]) );
DFFPOSX1 DFFPOSX1_1422 ( .CLK(clk_bF_buf85), .D(_282_), .Q(cpuregs_2_[0]) );
DFFPOSX1 DFFPOSX1_1423 ( .CLK(clk_bF_buf84), .D(_283_), .Q(cpuregs_2_[1]) );
DFFPOSX1 DFFPOSX1_1424 ( .CLK(clk_bF_buf83), .D(_284_), .Q(cpuregs_2_[2]) );
DFFPOSX1 DFFPOSX1_1425 ( .CLK(clk_bF_buf82), .D(_285_), .Q(cpuregs_2_[3]) );
DFFPOSX1 DFFPOSX1_1426 ( .CLK(clk_bF_buf81), .D(_286_), .Q(cpuregs_2_[4]) );
DFFPOSX1 DFFPOSX1_1427 ( .CLK(clk_bF_buf80), .D(_287_), .Q(cpuregs_2_[5]) );
DFFPOSX1 DFFPOSX1_1428 ( .CLK(clk_bF_buf79), .D(_288_), .Q(cpuregs_2_[6]) );
DFFPOSX1 DFFPOSX1_1429 ( .CLK(clk_bF_buf78), .D(_289_), .Q(cpuregs_2_[7]) );
DFFPOSX1 DFFPOSX1_1430 ( .CLK(clk_bF_buf77), .D(_290_), .Q(cpuregs_2_[8]) );
DFFPOSX1 DFFPOSX1_1431 ( .CLK(clk_bF_buf76), .D(_291_), .Q(cpuregs_2_[9]) );
DFFPOSX1 DFFPOSX1_1432 ( .CLK(clk_bF_buf75), .D(_292_), .Q(cpuregs_2_[10]) );
DFFPOSX1 DFFPOSX1_1433 ( .CLK(clk_bF_buf74), .D(_293_), .Q(cpuregs_2_[11]) );
DFFPOSX1 DFFPOSX1_1434 ( .CLK(clk_bF_buf73), .D(_294_), .Q(cpuregs_2_[12]) );
DFFPOSX1 DFFPOSX1_1435 ( .CLK(clk_bF_buf72), .D(_295_), .Q(cpuregs_2_[13]) );
DFFPOSX1 DFFPOSX1_1436 ( .CLK(clk_bF_buf71), .D(_296_), .Q(cpuregs_2_[14]) );
DFFPOSX1 DFFPOSX1_1437 ( .CLK(clk_bF_buf70), .D(_297_), .Q(cpuregs_2_[15]) );
DFFPOSX1 DFFPOSX1_1438 ( .CLK(clk_bF_buf69), .D(_298_), .Q(cpuregs_2_[16]) );
DFFPOSX1 DFFPOSX1_1439 ( .CLK(clk_bF_buf68), .D(_299_), .Q(cpuregs_2_[17]) );
DFFPOSX1 DFFPOSX1_1440 ( .CLK(clk_bF_buf67), .D(_300_), .Q(cpuregs_2_[18]) );
DFFPOSX1 DFFPOSX1_1441 ( .CLK(clk_bF_buf66), .D(_301_), .Q(cpuregs_2_[19]) );
DFFPOSX1 DFFPOSX1_1442 ( .CLK(clk_bF_buf65), .D(_302_), .Q(cpuregs_2_[20]) );
DFFPOSX1 DFFPOSX1_1443 ( .CLK(clk_bF_buf64), .D(_303_), .Q(cpuregs_2_[21]) );
DFFPOSX1 DFFPOSX1_1444 ( .CLK(clk_bF_buf63), .D(_304_), .Q(cpuregs_2_[22]) );
DFFPOSX1 DFFPOSX1_1445 ( .CLK(clk_bF_buf62), .D(_305_), .Q(cpuregs_2_[23]) );
DFFPOSX1 DFFPOSX1_1446 ( .CLK(clk_bF_buf61), .D(_306_), .Q(cpuregs_2_[24]) );
DFFPOSX1 DFFPOSX1_1447 ( .CLK(clk_bF_buf60), .D(_307_), .Q(cpuregs_2_[25]) );
DFFPOSX1 DFFPOSX1_1448 ( .CLK(clk_bF_buf59), .D(_308_), .Q(cpuregs_2_[26]) );
DFFPOSX1 DFFPOSX1_1449 ( .CLK(clk_bF_buf58), .D(_309_), .Q(cpuregs_2_[27]) );
DFFPOSX1 DFFPOSX1_1450 ( .CLK(clk_bF_buf57), .D(_310_), .Q(cpuregs_2_[28]) );
DFFPOSX1 DFFPOSX1_1451 ( .CLK(clk_bF_buf56), .D(_311_), .Q(cpuregs_2_[29]) );
DFFPOSX1 DFFPOSX1_1452 ( .CLK(clk_bF_buf55), .D(_312_), .Q(cpuregs_2_[30]) );
DFFPOSX1 DFFPOSX1_1453 ( .CLK(clk_bF_buf54), .D(_313_), .Q(cpuregs_2_[31]) );
DFFPOSX1 DFFPOSX1_1454 ( .CLK(clk_bF_buf53), .D(_122_), .Q(cpuregs_7_[0]) );
DFFPOSX1 DFFPOSX1_1455 ( .CLK(clk_bF_buf52), .D(_123_), .Q(cpuregs_7_[1]) );
DFFPOSX1 DFFPOSX1_1456 ( .CLK(clk_bF_buf51), .D(_124_), .Q(cpuregs_7_[2]) );
DFFPOSX1 DFFPOSX1_1457 ( .CLK(clk_bF_buf50), .D(_125_), .Q(cpuregs_7_[3]) );
DFFPOSX1 DFFPOSX1_1458 ( .CLK(clk_bF_buf49), .D(_126_), .Q(cpuregs_7_[4]) );
DFFPOSX1 DFFPOSX1_1459 ( .CLK(clk_bF_buf48), .D(_127_), .Q(cpuregs_7_[5]) );
DFFPOSX1 DFFPOSX1_1460 ( .CLK(clk_bF_buf47), .D(_128_), .Q(cpuregs_7_[6]) );
DFFPOSX1 DFFPOSX1_1461 ( .CLK(clk_bF_buf46), .D(_129_), .Q(cpuregs_7_[7]) );
DFFPOSX1 DFFPOSX1_1462 ( .CLK(clk_bF_buf45), .D(_130_), .Q(cpuregs_7_[8]) );
DFFPOSX1 DFFPOSX1_1463 ( .CLK(clk_bF_buf44), .D(_131_), .Q(cpuregs_7_[9]) );
DFFPOSX1 DFFPOSX1_1464 ( .CLK(clk_bF_buf43), .D(_132_), .Q(cpuregs_7_[10]) );
DFFPOSX1 DFFPOSX1_1465 ( .CLK(clk_bF_buf42), .D(_133_), .Q(cpuregs_7_[11]) );
DFFPOSX1 DFFPOSX1_1466 ( .CLK(clk_bF_buf41), .D(_134_), .Q(cpuregs_7_[12]) );
DFFPOSX1 DFFPOSX1_1467 ( .CLK(clk_bF_buf40), .D(_135_), .Q(cpuregs_7_[13]) );
DFFPOSX1 DFFPOSX1_1468 ( .CLK(clk_bF_buf39), .D(_136_), .Q(cpuregs_7_[14]) );
DFFPOSX1 DFFPOSX1_1469 ( .CLK(clk_bF_buf38), .D(_137_), .Q(cpuregs_7_[15]) );
DFFPOSX1 DFFPOSX1_1470 ( .CLK(clk_bF_buf37), .D(_138_), .Q(cpuregs_7_[16]) );
DFFPOSX1 DFFPOSX1_1471 ( .CLK(clk_bF_buf36), .D(_139_), .Q(cpuregs_7_[17]) );
DFFPOSX1 DFFPOSX1_1472 ( .CLK(clk_bF_buf35), .D(_140_), .Q(cpuregs_7_[18]) );
DFFPOSX1 DFFPOSX1_1473 ( .CLK(clk_bF_buf34), .D(_141_), .Q(cpuregs_7_[19]) );
DFFPOSX1 DFFPOSX1_1474 ( .CLK(clk_bF_buf33), .D(_142_), .Q(cpuregs_7_[20]) );
DFFPOSX1 DFFPOSX1_1475 ( .CLK(clk_bF_buf32), .D(_143_), .Q(cpuregs_7_[21]) );
DFFPOSX1 DFFPOSX1_1476 ( .CLK(clk_bF_buf31), .D(_144_), .Q(cpuregs_7_[22]) );
DFFPOSX1 DFFPOSX1_1477 ( .CLK(clk_bF_buf30), .D(_145_), .Q(cpuregs_7_[23]) );
DFFPOSX1 DFFPOSX1_1478 ( .CLK(clk_bF_buf29), .D(_146_), .Q(cpuregs_7_[24]) );
DFFPOSX1 DFFPOSX1_1479 ( .CLK(clk_bF_buf28), .D(_147_), .Q(cpuregs_7_[25]) );
DFFPOSX1 DFFPOSX1_1480 ( .CLK(clk_bF_buf27), .D(_148_), .Q(cpuregs_7_[26]) );
DFFPOSX1 DFFPOSX1_1481 ( .CLK(clk_bF_buf26), .D(_149_), .Q(cpuregs_7_[27]) );
DFFPOSX1 DFFPOSX1_1482 ( .CLK(clk_bF_buf25), .D(_150_), .Q(cpuregs_7_[28]) );
DFFPOSX1 DFFPOSX1_1483 ( .CLK(clk_bF_buf24), .D(_151_), .Q(cpuregs_7_[29]) );
DFFPOSX1 DFFPOSX1_1484 ( .CLK(clk_bF_buf23), .D(_152_), .Q(cpuregs_7_[30]) );
DFFPOSX1 DFFPOSX1_1485 ( .CLK(clk_bF_buf22), .D(_153_), .Q(cpuregs_7_[31]) );
DFFPOSX1 DFFPOSX1_1486 ( .CLK(clk_bF_buf21), .D(_250_), .Q(cpuregs_3_[0]) );
DFFPOSX1 DFFPOSX1_1487 ( .CLK(clk_bF_buf20), .D(_251_), .Q(cpuregs_3_[1]) );
DFFPOSX1 DFFPOSX1_1488 ( .CLK(clk_bF_buf19), .D(_252_), .Q(cpuregs_3_[2]) );
DFFPOSX1 DFFPOSX1_1489 ( .CLK(clk_bF_buf18), .D(_253_), .Q(cpuregs_3_[3]) );
DFFPOSX1 DFFPOSX1_1490 ( .CLK(clk_bF_buf17), .D(_254_), .Q(cpuregs_3_[4]) );
DFFPOSX1 DFFPOSX1_1491 ( .CLK(clk_bF_buf16), .D(_255_), .Q(cpuregs_3_[5]) );
DFFPOSX1 DFFPOSX1_1492 ( .CLK(clk_bF_buf15), .D(_256_), .Q(cpuregs_3_[6]) );
DFFPOSX1 DFFPOSX1_1493 ( .CLK(clk_bF_buf14), .D(_257_), .Q(cpuregs_3_[7]) );
DFFPOSX1 DFFPOSX1_1494 ( .CLK(clk_bF_buf13), .D(_258_), .Q(cpuregs_3_[8]) );
DFFPOSX1 DFFPOSX1_1495 ( .CLK(clk_bF_buf12), .D(_259_), .Q(cpuregs_3_[9]) );
DFFPOSX1 DFFPOSX1_1496 ( .CLK(clk_bF_buf11), .D(_260_), .Q(cpuregs_3_[10]) );
DFFPOSX1 DFFPOSX1_1497 ( .CLK(clk_bF_buf10), .D(_261_), .Q(cpuregs_3_[11]) );
DFFPOSX1 DFFPOSX1_1498 ( .CLK(clk_bF_buf9), .D(_262_), .Q(cpuregs_3_[12]) );
DFFPOSX1 DFFPOSX1_1499 ( .CLK(clk_bF_buf8), .D(_263_), .Q(cpuregs_3_[13]) );
DFFPOSX1 DFFPOSX1_1500 ( .CLK(clk_bF_buf7), .D(_264_), .Q(cpuregs_3_[14]) );
DFFPOSX1 DFFPOSX1_1501 ( .CLK(clk_bF_buf6), .D(_265_), .Q(cpuregs_3_[15]) );
DFFPOSX1 DFFPOSX1_1502 ( .CLK(clk_bF_buf5), .D(_266_), .Q(cpuregs_3_[16]) );
DFFPOSX1 DFFPOSX1_1503 ( .CLK(clk_bF_buf4), .D(_267_), .Q(cpuregs_3_[17]) );
DFFPOSX1 DFFPOSX1_1504 ( .CLK(clk_bF_buf3), .D(_268_), .Q(cpuregs_3_[18]) );
DFFPOSX1 DFFPOSX1_1505 ( .CLK(clk_bF_buf2), .D(_269_), .Q(cpuregs_3_[19]) );
DFFPOSX1 DFFPOSX1_1506 ( .CLK(clk_bF_buf1), .D(_270_), .Q(cpuregs_3_[20]) );
DFFPOSX1 DFFPOSX1_1507 ( .CLK(clk_bF_buf0), .D(_271_), .Q(cpuregs_3_[21]) );
DFFPOSX1 DFFPOSX1_1508 ( .CLK(clk_bF_buf136), .D(_272_), .Q(cpuregs_3_[22]) );
DFFPOSX1 DFFPOSX1_1509 ( .CLK(clk_bF_buf135), .D(_273_), .Q(cpuregs_3_[23]) );
DFFPOSX1 DFFPOSX1_1510 ( .CLK(clk_bF_buf134), .D(_274_), .Q(cpuregs_3_[24]) );
DFFPOSX1 DFFPOSX1_1511 ( .CLK(clk_bF_buf133), .D(_275_), .Q(cpuregs_3_[25]) );
DFFPOSX1 DFFPOSX1_1512 ( .CLK(clk_bF_buf132), .D(_276_), .Q(cpuregs_3_[26]) );
DFFPOSX1 DFFPOSX1_1513 ( .CLK(clk_bF_buf131), .D(_277_), .Q(cpuregs_3_[27]) );
DFFPOSX1 DFFPOSX1_1514 ( .CLK(clk_bF_buf130), .D(_278_), .Q(cpuregs_3_[28]) );
DFFPOSX1 DFFPOSX1_1515 ( .CLK(clk_bF_buf129), .D(_279_), .Q(cpuregs_3_[29]) );
DFFPOSX1 DFFPOSX1_1516 ( .CLK(clk_bF_buf128), .D(_280_), .Q(cpuregs_3_[30]) );
DFFPOSX1 DFFPOSX1_1517 ( .CLK(clk_bF_buf127), .D(_281_), .Q(cpuregs_3_[31]) );
DFFPOSX1 DFFPOSX1_1518 ( .CLK(clk_bF_buf126), .D(_1083_), .Q(cpuregs_13_[0]) );
DFFPOSX1 DFFPOSX1_1519 ( .CLK(clk_bF_buf125), .D(_1084_), .Q(cpuregs_13_[1]) );
DFFPOSX1 DFFPOSX1_1520 ( .CLK(clk_bF_buf124), .D(_1085_), .Q(cpuregs_13_[2]) );
DFFPOSX1 DFFPOSX1_1521 ( .CLK(clk_bF_buf123), .D(_1086_), .Q(cpuregs_13_[3]) );
DFFPOSX1 DFFPOSX1_1522 ( .CLK(clk_bF_buf122), .D(_1087_), .Q(cpuregs_13_[4]) );
DFFPOSX1 DFFPOSX1_1523 ( .CLK(clk_bF_buf121), .D(_1088_), .Q(cpuregs_13_[5]) );
DFFPOSX1 DFFPOSX1_1524 ( .CLK(clk_bF_buf120), .D(_1089_), .Q(cpuregs_13_[6]) );
DFFPOSX1 DFFPOSX1_1525 ( .CLK(clk_bF_buf119), .D(_1090_), .Q(cpuregs_13_[7]) );
DFFPOSX1 DFFPOSX1_1526 ( .CLK(clk_bF_buf118), .D(_1091_), .Q(cpuregs_13_[8]) );
DFFPOSX1 DFFPOSX1_1527 ( .CLK(clk_bF_buf117), .D(_1092_), .Q(cpuregs_13_[9]) );
DFFPOSX1 DFFPOSX1_1528 ( .CLK(clk_bF_buf116), .D(_1093_), .Q(cpuregs_13_[10]) );
DFFPOSX1 DFFPOSX1_1529 ( .CLK(clk_bF_buf115), .D(_1094_), .Q(cpuregs_13_[11]) );
DFFPOSX1 DFFPOSX1_1530 ( .CLK(clk_bF_buf114), .D(_1095_), .Q(cpuregs_13_[12]) );
DFFPOSX1 DFFPOSX1_1531 ( .CLK(clk_bF_buf113), .D(_1096_), .Q(cpuregs_13_[13]) );
DFFPOSX1 DFFPOSX1_1532 ( .CLK(clk_bF_buf112), .D(_1097_), .Q(cpuregs_13_[14]) );
DFFPOSX1 DFFPOSX1_1533 ( .CLK(clk_bF_buf111), .D(_1098_), .Q(cpuregs_13_[15]) );
DFFPOSX1 DFFPOSX1_1534 ( .CLK(clk_bF_buf110), .D(_1099_), .Q(cpuregs_13_[16]) );
DFFPOSX1 DFFPOSX1_1535 ( .CLK(clk_bF_buf109), .D(_1100_), .Q(cpuregs_13_[17]) );
DFFPOSX1 DFFPOSX1_1536 ( .CLK(clk_bF_buf108), .D(_1101_), .Q(cpuregs_13_[18]) );
DFFPOSX1 DFFPOSX1_1537 ( .CLK(clk_bF_buf107), .D(_1102_), .Q(cpuregs_13_[19]) );
DFFPOSX1 DFFPOSX1_1538 ( .CLK(clk_bF_buf106), .D(_1103_), .Q(cpuregs_13_[20]) );
DFFPOSX1 DFFPOSX1_1539 ( .CLK(clk_bF_buf105), .D(_1104_), .Q(cpuregs_13_[21]) );
DFFPOSX1 DFFPOSX1_1540 ( .CLK(clk_bF_buf104), .D(_1105_), .Q(cpuregs_13_[22]) );
DFFPOSX1 DFFPOSX1_1541 ( .CLK(clk_bF_buf103), .D(_1106_), .Q(cpuregs_13_[23]) );
DFFPOSX1 DFFPOSX1_1542 ( .CLK(clk_bF_buf102), .D(_1107_), .Q(cpuregs_13_[24]) );
DFFPOSX1 DFFPOSX1_1543 ( .CLK(clk_bF_buf101), .D(_1108_), .Q(cpuregs_13_[25]) );
DFFPOSX1 DFFPOSX1_1544 ( .CLK(clk_bF_buf100), .D(_1109_), .Q(cpuregs_13_[26]) );
DFFPOSX1 DFFPOSX1_1545 ( .CLK(clk_bF_buf99), .D(_1110_), .Q(cpuregs_13_[27]) );
DFFPOSX1 DFFPOSX1_1546 ( .CLK(clk_bF_buf98), .D(_1111_), .Q(cpuregs_13_[28]) );
DFFPOSX1 DFFPOSX1_1547 ( .CLK(clk_bF_buf97), .D(_1112_), .Q(cpuregs_13_[29]) );
DFFPOSX1 DFFPOSX1_1548 ( .CLK(clk_bF_buf96), .D(_1113_), .Q(cpuregs_13_[30]) );
DFFPOSX1 DFFPOSX1_1549 ( .CLK(clk_bF_buf95), .D(_1114_), .Q(cpuregs_13_[31]) );
DFFPOSX1 DFFPOSX1_1550 ( .CLK(clk_bF_buf94), .D(_731_), .Q(cpuregs_10_[0]) );
DFFPOSX1 DFFPOSX1_1551 ( .CLK(clk_bF_buf93), .D(_732_), .Q(cpuregs_10_[1]) );
DFFPOSX1 DFFPOSX1_1552 ( .CLK(clk_bF_buf92), .D(_733_), .Q(cpuregs_10_[2]) );
DFFPOSX1 DFFPOSX1_1553 ( .CLK(clk_bF_buf91), .D(_734_), .Q(cpuregs_10_[3]) );
DFFPOSX1 DFFPOSX1_1554 ( .CLK(clk_bF_buf90), .D(_735_), .Q(cpuregs_10_[4]) );
DFFPOSX1 DFFPOSX1_1555 ( .CLK(clk_bF_buf89), .D(_736_), .Q(cpuregs_10_[5]) );
DFFPOSX1 DFFPOSX1_1556 ( .CLK(clk_bF_buf88), .D(_737_), .Q(cpuregs_10_[6]) );
DFFPOSX1 DFFPOSX1_1557 ( .CLK(clk_bF_buf87), .D(_738_), .Q(cpuregs_10_[7]) );
DFFPOSX1 DFFPOSX1_1558 ( .CLK(clk_bF_buf86), .D(_739_), .Q(cpuregs_10_[8]) );
DFFPOSX1 DFFPOSX1_1559 ( .CLK(clk_bF_buf85), .D(_740_), .Q(cpuregs_10_[9]) );
DFFPOSX1 DFFPOSX1_1560 ( .CLK(clk_bF_buf84), .D(_741_), .Q(cpuregs_10_[10]) );
DFFPOSX1 DFFPOSX1_1561 ( .CLK(clk_bF_buf83), .D(_742_), .Q(cpuregs_10_[11]) );
DFFPOSX1 DFFPOSX1_1562 ( .CLK(clk_bF_buf82), .D(_743_), .Q(cpuregs_10_[12]) );
DFFPOSX1 DFFPOSX1_1563 ( .CLK(clk_bF_buf81), .D(_744_), .Q(cpuregs_10_[13]) );
DFFPOSX1 DFFPOSX1_1564 ( .CLK(clk_bF_buf80), .D(_745_), .Q(cpuregs_10_[14]) );
DFFPOSX1 DFFPOSX1_1565 ( .CLK(clk_bF_buf79), .D(_746_), .Q(cpuregs_10_[15]) );
DFFPOSX1 DFFPOSX1_1566 ( .CLK(clk_bF_buf78), .D(_747_), .Q(cpuregs_10_[16]) );
DFFPOSX1 DFFPOSX1_1567 ( .CLK(clk_bF_buf77), .D(_748_), .Q(cpuregs_10_[17]) );
DFFPOSX1 DFFPOSX1_1568 ( .CLK(clk_bF_buf76), .D(_749_), .Q(cpuregs_10_[18]) );
DFFPOSX1 DFFPOSX1_1569 ( .CLK(clk_bF_buf75), .D(_750_), .Q(cpuregs_10_[19]) );
DFFPOSX1 DFFPOSX1_1570 ( .CLK(clk_bF_buf74), .D(_751_), .Q(cpuregs_10_[20]) );
DFFPOSX1 DFFPOSX1_1571 ( .CLK(clk_bF_buf73), .D(_752_), .Q(cpuregs_10_[21]) );
DFFPOSX1 DFFPOSX1_1572 ( .CLK(clk_bF_buf72), .D(_753_), .Q(cpuregs_10_[22]) );
DFFPOSX1 DFFPOSX1_1573 ( .CLK(clk_bF_buf71), .D(_754_), .Q(cpuregs_10_[23]) );
DFFPOSX1 DFFPOSX1_1574 ( .CLK(clk_bF_buf70), .D(_755_), .Q(cpuregs_10_[24]) );
DFFPOSX1 DFFPOSX1_1575 ( .CLK(clk_bF_buf69), .D(_756_), .Q(cpuregs_10_[25]) );
DFFPOSX1 DFFPOSX1_1576 ( .CLK(clk_bF_buf68), .D(_757_), .Q(cpuregs_10_[26]) );
DFFPOSX1 DFFPOSX1_1577 ( .CLK(clk_bF_buf67), .D(_758_), .Q(cpuregs_10_[27]) );
DFFPOSX1 DFFPOSX1_1578 ( .CLK(clk_bF_buf66), .D(_759_), .Q(cpuregs_10_[28]) );
DFFPOSX1 DFFPOSX1_1579 ( .CLK(clk_bF_buf65), .D(_760_), .Q(cpuregs_10_[29]) );
DFFPOSX1 DFFPOSX1_1580 ( .CLK(clk_bF_buf64), .D(_761_), .Q(cpuregs_10_[30]) );
DFFPOSX1 DFFPOSX1_1581 ( .CLK(clk_bF_buf63), .D(_762_), .Q(cpuregs_10_[31]) );
DFFPOSX1 DFFPOSX1_1582 ( .CLK(clk_bF_buf62), .D(_667_), .Q(cpuregs_22_[0]) );
DFFPOSX1 DFFPOSX1_1583 ( .CLK(clk_bF_buf61), .D(_668_), .Q(cpuregs_22_[1]) );
DFFPOSX1 DFFPOSX1_1584 ( .CLK(clk_bF_buf60), .D(_669_), .Q(cpuregs_22_[2]) );
DFFPOSX1 DFFPOSX1_1585 ( .CLK(clk_bF_buf59), .D(_670_), .Q(cpuregs_22_[3]) );
DFFPOSX1 DFFPOSX1_1586 ( .CLK(clk_bF_buf58), .D(_671_), .Q(cpuregs_22_[4]) );
DFFPOSX1 DFFPOSX1_1587 ( .CLK(clk_bF_buf57), .D(_672_), .Q(cpuregs_22_[5]) );
DFFPOSX1 DFFPOSX1_1588 ( .CLK(clk_bF_buf56), .D(_673_), .Q(cpuregs_22_[6]) );
DFFPOSX1 DFFPOSX1_1589 ( .CLK(clk_bF_buf55), .D(_674_), .Q(cpuregs_22_[7]) );
DFFPOSX1 DFFPOSX1_1590 ( .CLK(clk_bF_buf54), .D(_675_), .Q(cpuregs_22_[8]) );
DFFPOSX1 DFFPOSX1_1591 ( .CLK(clk_bF_buf53), .D(_676_), .Q(cpuregs_22_[9]) );
DFFPOSX1 DFFPOSX1_1592 ( .CLK(clk_bF_buf52), .D(_677_), .Q(cpuregs_22_[10]) );
DFFPOSX1 DFFPOSX1_1593 ( .CLK(clk_bF_buf51), .D(_678_), .Q(cpuregs_22_[11]) );
DFFPOSX1 DFFPOSX1_1594 ( .CLK(clk_bF_buf50), .D(_679_), .Q(cpuregs_22_[12]) );
DFFPOSX1 DFFPOSX1_1595 ( .CLK(clk_bF_buf49), .D(_680_), .Q(cpuregs_22_[13]) );
DFFPOSX1 DFFPOSX1_1596 ( .CLK(clk_bF_buf48), .D(_681_), .Q(cpuregs_22_[14]) );
DFFPOSX1 DFFPOSX1_1597 ( .CLK(clk_bF_buf47), .D(_682_), .Q(cpuregs_22_[15]) );
DFFPOSX1 DFFPOSX1_1598 ( .CLK(clk_bF_buf46), .D(_683_), .Q(cpuregs_22_[16]) );
DFFPOSX1 DFFPOSX1_1599 ( .CLK(clk_bF_buf45), .D(_684_), .Q(cpuregs_22_[17]) );
DFFPOSX1 DFFPOSX1_1600 ( .CLK(clk_bF_buf44), .D(_685_), .Q(cpuregs_22_[18]) );
DFFPOSX1 DFFPOSX1_1601 ( .CLK(clk_bF_buf43), .D(_686_), .Q(cpuregs_22_[19]) );
DFFPOSX1 DFFPOSX1_1602 ( .CLK(clk_bF_buf42), .D(_687_), .Q(cpuregs_22_[20]) );
DFFPOSX1 DFFPOSX1_1603 ( .CLK(clk_bF_buf41), .D(_688_), .Q(cpuregs_22_[21]) );
DFFPOSX1 DFFPOSX1_1604 ( .CLK(clk_bF_buf40), .D(_689_), .Q(cpuregs_22_[22]) );
DFFPOSX1 DFFPOSX1_1605 ( .CLK(clk_bF_buf39), .D(_690_), .Q(cpuregs_22_[23]) );
DFFPOSX1 DFFPOSX1_1606 ( .CLK(clk_bF_buf38), .D(_691_), .Q(cpuregs_22_[24]) );
DFFPOSX1 DFFPOSX1_1607 ( .CLK(clk_bF_buf37), .D(_692_), .Q(cpuregs_22_[25]) );
DFFPOSX1 DFFPOSX1_1608 ( .CLK(clk_bF_buf36), .D(_693_), .Q(cpuregs_22_[26]) );
DFFPOSX1 DFFPOSX1_1609 ( .CLK(clk_bF_buf35), .D(_694_), .Q(cpuregs_22_[27]) );
DFFPOSX1 DFFPOSX1_1610 ( .CLK(clk_bF_buf34), .D(_695_), .Q(cpuregs_22_[28]) );
DFFPOSX1 DFFPOSX1_1611 ( .CLK(clk_bF_buf33), .D(_696_), .Q(cpuregs_22_[29]) );
DFFPOSX1 DFFPOSX1_1612 ( .CLK(clk_bF_buf32), .D(_697_), .Q(cpuregs_22_[30]) );
DFFPOSX1 DFFPOSX1_1613 ( .CLK(clk_bF_buf31), .D(_698_), .Q(cpuregs_22_[31]) );
endmodule
